module database#(
parameter maxl=5,
parameter sizein=40,
parameter sizew=8
)
(
input clk,
input rst,

input[7:0] rnum,//the number
input[7:0] rsam,//the sample
input[7:0] rlayer,//the layer to be read
input[7:0] rn,//the neuron to be read
input[7:0] rin,//the input of a neuron
input rmode,//0: read input, 1: read weight/bias
input rs,//start
output reg[sizein-1:0] ram_in,
output reg[sizew-1:0] ram_w,
output reg rf//finished
);

parameter IDLE=0;
parameter ADDR=1;
parameter WAIT=2;
parameter READ=3;

reg [7:0] state;

always@(posedge clk)begin
	if(rst)begin
		ram_in<=0;
		ram_w<=0;
		rf<=0;
		state<=IDLE;
	end
	else begin
		case(state)
		IDLE:begin
			if(rs)begin
				ram_in<=0;
				ram_w<=0;
				rf<=0;
				state<=WAIT;
			end
			else begin
				state<=IDLE;
			end
		end
		WAIT:begin
			state<=READ;
		end
		READ:begin
			if(rmode==0)begin
				case({rnum,rsam,rin})
0:begin
	ram_in<=32'd256;
end
1:begin
	ram_in<=32'd896;
end
2:begin
	ram_in<=32'd960;
end
3:begin
	ram_in<=32'd1984;
end
4:begin
	ram_in<=32'd4064;
end
5:begin
	ram_in<=32'd3936;
end
6:begin
	ram_in<=32'd3616;
end
7:begin
	ram_in<=32'd3616;
end
8:begin
	ram_in<=32'd7200;
end
9:begin
	ram_in<=32'd7216;
end
10:begin
	ram_in<=32'd7184;
end
11:begin
	ram_in<=32'd7184;
end
12:begin
	ram_in<=32'd7192;
end
13:begin
	ram_in<=32'd7192;
end
14:begin
	ram_in<=32'd3080;
end
15:begin
	ram_in<=32'd3080;
end
16:begin
	ram_in<=32'd3080;
end
17:begin
	ram_in<=32'd7176;
end
18:begin
	ram_in<=32'd7176;
end
19:begin
	ram_in<=32'd3084;
end
20:begin
	ram_in<=32'd3084;
end
21:begin
	ram_in<=32'd3084;
end
22:begin
	ram_in<=32'd3100;
end
23:begin
	ram_in<=32'd1548;
end
24:begin
	ram_in<=32'd1564;
end
25:begin
	ram_in<=32'd1564;
end
26:begin
	ram_in<=32'd1592;
end
27:begin
	ram_in<=32'd1912;
end
28:begin
	ram_in<=32'd1016;
end
29:begin
	ram_in<=32'd1008;
end
30:begin
	ram_in<=32'd992;
end
31:begin
	ram_in<=32'd448;
end
256:begin
	ram_in<=32'd128;
end
257:begin
	ram_in<=32'd960;
end
258:begin
	ram_in<=32'd2016;
end
259:begin
	ram_in<=32'd2016;
end
260:begin
	ram_in<=32'd2032;
end
261:begin
	ram_in<=32'd1904;
end
262:begin
	ram_in<=32'd3632;
end
263:begin
	ram_in<=32'd3632;
end
264:begin
	ram_in<=32'd3640;
end
265:begin
	ram_in<=32'd3640;
end
266:begin
	ram_in<=32'd3608;
end
267:begin
	ram_in<=32'd3608;
end
268:begin
	ram_in<=32'd3612;
end
269:begin
	ram_in<=32'd3096;
end
270:begin
	ram_in<=32'd3096;
end
271:begin
	ram_in<=32'd3096;
end
272:begin
	ram_in<=32'd3080;
end
273:begin
	ram_in<=32'd3080;
end
274:begin
	ram_in<=32'd3080;
end
275:begin
	ram_in<=32'd3080;
end
276:begin
	ram_in<=32'd3096;
end
277:begin
	ram_in<=32'd3096;
end
278:begin
	ram_in<=32'd3096;
end
279:begin
	ram_in<=32'd3704;
end
280:begin
	ram_in<=32'd3824;
end
281:begin
	ram_in<=32'd4080;
end
282:begin
	ram_in<=32'd2032;
end
283:begin
	ram_in<=32'd4064;
end
284:begin
	ram_in<=32'd1984;
end
285:begin
	ram_in<=32'd1920;
end
286:begin
	ram_in<=32'd1792;
end
287:begin
	ram_in<=32'd0;
end
512:begin
	ram_in<=32'd512;
end
513:begin
	ram_in<=32'd1536;
end
514:begin
	ram_in<=32'd1920;
end
515:begin
	ram_in<=32'd1984;
end
516:begin
	ram_in<=32'd1984;
end
517:begin
	ram_in<=32'd4064;
end
518:begin
	ram_in<=32'd4064;
end
519:begin
	ram_in<=32'd3936;
end
520:begin
	ram_in<=32'd3680;
end
521:begin
	ram_in<=32'd3632;
end
522:begin
	ram_in<=32'd3608;
end
523:begin
	ram_in<=32'd3608;
end
524:begin
	ram_in<=32'd3608;
end
525:begin
	ram_in<=32'd3608;
end
526:begin
	ram_in<=32'd3096;
end
527:begin
	ram_in<=32'd3080;
end
528:begin
	ram_in<=32'd7176;
end
529:begin
	ram_in<=32'd7176;
end
530:begin
	ram_in<=32'd6168;
end
531:begin
	ram_in<=32'd6168;
end
532:begin
	ram_in<=32'd6168;
end
533:begin
	ram_in<=32'd6168;
end
534:begin
	ram_in<=32'd2072;
end
535:begin
	ram_in<=32'd3096;
end
536:begin
	ram_in<=32'd3128;
end
537:begin
	ram_in<=32'd3184;
end
538:begin
	ram_in<=32'd3184;
end
539:begin
	ram_in<=32'd4080;
end
540:begin
	ram_in<=32'd2016;
end
541:begin
	ram_in<=32'd1984;
end
542:begin
	ram_in<=32'd1984;
end
543:begin
	ram_in<=32'd768;
end
768:begin
	ram_in<=32'd256;
end
769:begin
	ram_in<=32'd384;
end
770:begin
	ram_in<=32'd896;
end
771:begin
	ram_in<=32'd960;
end
772:begin
	ram_in<=32'd1984;
end
773:begin
	ram_in<=32'd1888;
end
774:begin
	ram_in<=32'd1632;
end
775:begin
	ram_in<=32'd3680;
end
776:begin
	ram_in<=32'd3616;
end
777:begin
	ram_in<=32'd3632;
end
778:begin
	ram_in<=32'd3632;
end
779:begin
	ram_in<=32'd3608;
end
780:begin
	ram_in<=32'd3096;
end
781:begin
	ram_in<=32'd3096;
end
782:begin
	ram_in<=32'd3096;
end
783:begin
	ram_in<=32'd3592;
end
784:begin
	ram_in<=32'd3080;
end
785:begin
	ram_in<=32'd3080;
end
786:begin
	ram_in<=32'd3596;
end
787:begin
	ram_in<=32'd3596;
end
788:begin
	ram_in<=32'd3596;
end
789:begin
	ram_in<=32'd3612;
end
790:begin
	ram_in<=32'd1820;
end
791:begin
	ram_in<=32'd1820;
end
792:begin
	ram_in<=32'd1080;
end
793:begin
	ram_in<=32'd1592;
end
794:begin
	ram_in<=32'd1656;
end
795:begin
	ram_in<=32'd2032;
end
796:begin
	ram_in<=32'd1008;
end
797:begin
	ram_in<=32'd992;
end
798:begin
	ram_in<=32'd960;
end
799:begin
	ram_in<=32'd256;
end
1024:begin
	ram_in<=32'd384;
end
1025:begin
	ram_in<=32'd992;
end
1026:begin
	ram_in<=32'd1760;
end
1027:begin
	ram_in<=32'd1776;
end
1028:begin
	ram_in<=32'd4080;
end
1029:begin
	ram_in<=32'd4080;
end
1030:begin
	ram_in<=32'd3632;
end
1031:begin
	ram_in<=32'd7216;
end
1032:begin
	ram_in<=32'd7192;
end
1033:begin
	ram_in<=32'd7192;
end
1034:begin
	ram_in<=32'd7688;
end
1035:begin
	ram_in<=32'd7688;
end
1036:begin
	ram_in<=32'd7176;
end
1037:begin
	ram_in<=32'd7176;
end
1038:begin
	ram_in<=32'd3096;
end
1039:begin
	ram_in<=32'd3096;
end
1040:begin
	ram_in<=32'd3096;
end
1041:begin
	ram_in<=32'd3096;
end
1042:begin
	ram_in<=32'd3096;
end
1043:begin
	ram_in<=32'd2072;
end
1044:begin
	ram_in<=32'd2072;
end
1045:begin
	ram_in<=32'd2096;
end
1046:begin
	ram_in<=32'd6192;
end
1047:begin
	ram_in<=32'd3128;
end
1048:begin
	ram_in<=32'd3120;
end
1049:begin
	ram_in<=32'd3184;
end
1050:begin
	ram_in<=32'd3696;
end
1051:begin
	ram_in<=32'd2032;
end
1052:begin
	ram_in<=32'd2016;
end
1053:begin
	ram_in<=32'd1984;
end
1054:begin
	ram_in<=32'd1984;
end
1055:begin
	ram_in<=32'd384;
end
1280:begin
	ram_in<=32'd256;
end
1281:begin
	ram_in<=32'd896;
end
1282:begin
	ram_in<=32'd960;
end
1283:begin
	ram_in<=32'd1984;
end
1284:begin
	ram_in<=32'd4064;
end
1285:begin
	ram_in<=32'd4064;
end
1286:begin
	ram_in<=32'd4080;
end
1287:begin
	ram_in<=32'd3888;
end
1288:begin
	ram_in<=32'd3632;
end
1289:begin
	ram_in<=32'd7216;
end
1290:begin
	ram_in<=32'd7224;
end
1291:begin
	ram_in<=32'd7192;
end
1292:begin
	ram_in<=32'd7192;
end
1293:begin
	ram_in<=32'd3608;
end
1294:begin
	ram_in<=32'd7704;
end
1295:begin
	ram_in<=32'd7192;
end
1296:begin
	ram_in<=32'd3096;
end
1297:begin
	ram_in<=32'd7192;
end
1298:begin
	ram_in<=32'd3096;
end
1299:begin
	ram_in<=32'd3096;
end
1300:begin
	ram_in<=32'd3612;
end
1301:begin
	ram_in<=32'd3612;
end
1302:begin
	ram_in<=32'd3612;
end
1303:begin
	ram_in<=32'd3608;
end
1304:begin
	ram_in<=32'd3640;
end
1305:begin
	ram_in<=32'd3640;
end
1306:begin
	ram_in<=32'd2040;
end
1307:begin
	ram_in<=32'd2040;
end
1308:begin
	ram_in<=32'd2040;
end
1309:begin
	ram_in<=32'd1008;
end
1310:begin
	ram_in<=32'd992;
end
1311:begin
	ram_in<=32'd448;
end
1536:begin
	ram_in<=32'd0;
end
1537:begin
	ram_in<=32'd448;
end
1538:begin
	ram_in<=32'd960;
end
1539:begin
	ram_in<=32'd992;
end
1540:begin
	ram_in<=32'd2016;
end
1541:begin
	ram_in<=32'd2032;
end
1542:begin
	ram_in<=32'd3952;
end
1543:begin
	ram_in<=32'd3632;
end
1544:begin
	ram_in<=32'd3632;
end
1545:begin
	ram_in<=32'd7184;
end
1546:begin
	ram_in<=32'd6160;
end
1547:begin
	ram_in<=32'd7192;
end
1548:begin
	ram_in<=32'd6168;
end
1549:begin
	ram_in<=32'd6168;
end
1550:begin
	ram_in<=32'd6168;
end
1551:begin
	ram_in<=32'd3080;
end
1552:begin
	ram_in<=32'd6168;
end
1553:begin
	ram_in<=32'd6168;
end
1554:begin
	ram_in<=32'd3080;
end
1555:begin
	ram_in<=32'd3096;
end
1556:begin
	ram_in<=32'd3096;
end
1557:begin
	ram_in<=32'd3096;
end
1558:begin
	ram_in<=32'd3096;
end
1559:begin
	ram_in<=32'd1048;
end
1560:begin
	ram_in<=32'd1592;
end
1561:begin
	ram_in<=32'd1592;
end
1562:begin
	ram_in<=32'd1848;
end
1563:begin
	ram_in<=32'd2032;
end
1564:begin
	ram_in<=32'd1008;
end
1565:begin
	ram_in<=32'd1008;
end
1566:begin
	ram_in<=32'd496;
end
1567:begin
	ram_in<=32'd64;
end
1792:begin
	ram_in<=32'd384;
end
1793:begin
	ram_in<=32'd960;
end
1794:begin
	ram_in<=32'd1984;
end
1795:begin
	ram_in<=32'd1984;
end
1796:begin
	ram_in<=32'd2016;
end
1797:begin
	ram_in<=32'd2032;
end
1798:begin
	ram_in<=32'd2032;
end
1799:begin
	ram_in<=32'd4080;
end
1800:begin
	ram_in<=32'd4088;
end
1801:begin
	ram_in<=32'd4024;
end
1802:begin
	ram_in<=32'd3992;
end
1803:begin
	ram_in<=32'd3864;
end
1804:begin
	ram_in<=32'd6936;
end
1805:begin
	ram_in<=32'd3336;
end
1806:begin
	ram_in<=32'd3336;
end
1807:begin
	ram_in<=32'd3080;
end
1808:begin
	ram_in<=32'd6152;
end
1809:begin
	ram_in<=32'd6168;
end
1810:begin
	ram_in<=32'd6168;
end
1811:begin
	ram_in<=32'd6168;
end
1812:begin
	ram_in<=32'd3100;
end
1813:begin
	ram_in<=32'd3096;
end
1814:begin
	ram_in<=32'd3096;
end
1815:begin
	ram_in<=32'd3128;
end
1816:begin
	ram_in<=32'd3128;
end
1817:begin
	ram_in<=32'd3184;
end
1818:begin
	ram_in<=32'd4080;
end
1819:begin
	ram_in<=32'd2032;
end
1820:begin
	ram_in<=32'd2016;
end
1821:begin
	ram_in<=32'd2016;
end
1822:begin
	ram_in<=32'd960;
end
1823:begin
	ram_in<=32'd384;
end
2048:begin
	ram_in<=32'd256;
end
2049:begin
	ram_in<=32'd896;
end
2050:begin
	ram_in<=32'd1920;
end
2051:begin
	ram_in<=32'd1920;
end
2052:begin
	ram_in<=32'd1920;
end
2053:begin
	ram_in<=32'd2016;
end
2054:begin
	ram_in<=32'd2032;
end
2055:begin
	ram_in<=32'd2032;
end
2056:begin
	ram_in<=32'd4080;
end
2057:begin
	ram_in<=32'd4088;
end
2058:begin
	ram_in<=32'd4088;
end
2059:begin
	ram_in<=32'd3896;
end
2060:begin
	ram_in<=32'd3608;
end
2061:begin
	ram_in<=32'd3080;
end
2062:begin
	ram_in<=32'd3080;
end
2063:begin
	ram_in<=32'd3080;
end
2064:begin
	ram_in<=32'd2056;
end
2065:begin
	ram_in<=32'd2056;
end
2066:begin
	ram_in<=32'd6152;
end
2067:begin
	ram_in<=32'd6152;
end
2068:begin
	ram_in<=32'd3084;
end
2069:begin
	ram_in<=32'd3100;
end
2070:begin
	ram_in<=32'd3100;
end
2071:begin
	ram_in<=32'd3132;
end
2072:begin
	ram_in<=32'd3128;
end
2073:begin
	ram_in<=32'd3832;
end
2074:begin
	ram_in<=32'd4088;
end
2075:begin
	ram_in<=32'd2040;
end
2076:begin
	ram_in<=32'd2032;
end
2077:begin
	ram_in<=32'd2032;
end
2078:begin
	ram_in<=32'd992;
end
2079:begin
	ram_in<=32'd896;
end
2304:begin
	ram_in<=32'd512;
end
2305:begin
	ram_in<=32'd512;
end
2306:begin
	ram_in<=32'd1984;
end
2307:begin
	ram_in<=32'd2016;
end
2308:begin
	ram_in<=32'd2016;
end
2309:begin
	ram_in<=32'd4080;
end
2310:begin
	ram_in<=32'd4080;
end
2311:begin
	ram_in<=32'd4080;
end
2312:begin
	ram_in<=32'd3856;
end
2313:begin
	ram_in<=32'd3608;
end
2314:begin
	ram_in<=32'd3608;
end
2315:begin
	ram_in<=32'd3608;
end
2316:begin
	ram_in<=32'd2056;
end
2317:begin
	ram_in<=32'd2056;
end
2318:begin
	ram_in<=32'd2056;
end
2319:begin
	ram_in<=32'd2056;
end
2320:begin
	ram_in<=32'd6152;
end
2321:begin
	ram_in<=32'd6152;
end
2322:begin
	ram_in<=32'd6152;
end
2323:begin
	ram_in<=32'd6168;
end
2324:begin
	ram_in<=32'd6168;
end
2325:begin
	ram_in<=32'd2072;
end
2326:begin
	ram_in<=32'd2072;
end
2327:begin
	ram_in<=32'd2104;
end
2328:begin
	ram_in<=32'd3192;
end
2329:begin
	ram_in<=32'd3184;
end
2330:begin
	ram_in<=32'd3312;
end
2331:begin
	ram_in<=32'd4064;
end
2332:begin
	ram_in<=32'd1984;
end
2333:begin
	ram_in<=32'd1984;
end
2334:begin
	ram_in<=32'd960;
end
2335:begin
	ram_in<=32'd768;
end
65536:begin
	ram_in<=32'd0;
end
65537:begin
	ram_in<=32'd896;
end
65538:begin
	ram_in<=32'd992;
end
65539:begin
	ram_in<=32'd992;
end
65540:begin
	ram_in<=32'd992;
end
65541:begin
	ram_in<=32'd992;
end
65542:begin
	ram_in<=32'd2016;
end
65543:begin
	ram_in<=32'd2016;
end
65544:begin
	ram_in<=32'd1984;
end
65545:begin
	ram_in<=32'd1984;
end
65546:begin
	ram_in<=32'd1984;
end
65547:begin
	ram_in<=32'd1984;
end
65548:begin
	ram_in<=32'd2016;
end
65549:begin
	ram_in<=32'd4032;
end
65550:begin
	ram_in<=32'd4032;
end
65551:begin
	ram_in<=32'd4032;
end
65552:begin
	ram_in<=32'd8128;
end
65553:begin
	ram_in<=32'd8128;
end
65554:begin
	ram_in<=32'd4032;
end
65555:begin
	ram_in<=32'd4032;
end
65556:begin
	ram_in<=32'd3968;
end
65557:begin
	ram_in<=32'd1984;
end
65558:begin
	ram_in<=32'd1920;
end
65559:begin
	ram_in<=32'd1984;
end
65560:begin
	ram_in<=32'd1984;
end
65561:begin
	ram_in<=32'd1984;
end
65562:begin
	ram_in<=32'd1984;
end
65563:begin
	ram_in<=32'd960;
end
65564:begin
	ram_in<=32'd2016;
end
65565:begin
	ram_in<=32'd1008;
end
65566:begin
	ram_in<=32'd1008;
end
65567:begin
	ram_in<=32'd496;
end
65792:begin
	ram_in<=32'd224;
end
65793:begin
	ram_in<=32'd224;
end
65794:begin
	ram_in<=32'd240;
end
65795:begin
	ram_in<=32'd240;
end
65796:begin
	ram_in<=32'd496;
end
65797:begin
	ram_in<=32'd240;
end
65798:begin
	ram_in<=32'd240;
end
65799:begin
	ram_in<=32'd480;
end
65800:begin
	ram_in<=32'd480;
end
65801:begin
	ram_in<=32'd480;
end
65802:begin
	ram_in<=32'd480;
end
65803:begin
	ram_in<=32'd480;
end
65804:begin
	ram_in<=32'd480;
end
65805:begin
	ram_in<=32'd960;
end
65806:begin
	ram_in<=32'd1984;
end
65807:begin
	ram_in<=32'd4032;
end
65808:begin
	ram_in<=32'd8128;
end
65809:begin
	ram_in<=32'd8128;
end
65810:begin
	ram_in<=32'd8128;
end
65811:begin
	ram_in<=32'd1984;
end
65812:begin
	ram_in<=32'd448;
end
65813:begin
	ram_in<=32'd448;
end
65814:begin
	ram_in<=32'd960;
end
65815:begin
	ram_in<=32'd960;
end
65816:begin
	ram_in<=32'd960;
end
65817:begin
	ram_in<=32'd992;
end
65818:begin
	ram_in<=32'd992;
end
65819:begin
	ram_in<=32'd480;
end
65820:begin
	ram_in<=32'd248;
end
65821:begin
	ram_in<=32'd248;
end
65822:begin
	ram_in<=32'd120;
end
65823:begin
	ram_in<=32'd48;
end
66048:begin
	ram_in<=32'd768;
end
66049:begin
	ram_in<=32'd960;
end
66050:begin
	ram_in<=32'd992;
end
66051:begin
	ram_in<=32'd992;
end
66052:begin
	ram_in<=32'd480;
end
66053:begin
	ram_in<=32'd992;
end
66054:begin
	ram_in<=32'd2016;
end
66055:begin
	ram_in<=32'd992;
end
66056:begin
	ram_in<=32'd1984;
end
66057:begin
	ram_in<=32'd1984;
end
66058:begin
	ram_in<=32'd1984;
end
66059:begin
	ram_in<=32'd1984;
end
66060:begin
	ram_in<=32'd1984;
end
66061:begin
	ram_in<=32'd1984;
end
66062:begin
	ram_in<=32'd3968;
end
66063:begin
	ram_in<=32'd4032;
end
66064:begin
	ram_in<=32'd4032;
end
66065:begin
	ram_in<=32'd8064;
end
66066:begin
	ram_in<=32'd4032;
end
66067:begin
	ram_in<=32'd4032;
end
66068:begin
	ram_in<=32'd3968;
end
66069:begin
	ram_in<=32'd1792;
end
66070:begin
	ram_in<=32'd1984;
end
66071:begin
	ram_in<=32'd960;
end
66072:begin
	ram_in<=32'd960;
end
66073:begin
	ram_in<=32'd896;
end
66074:begin
	ram_in<=32'd960;
end
66075:begin
	ram_in<=32'd992;
end
66076:begin
	ram_in<=32'd992;
end
66077:begin
	ram_in<=32'd992;
end
66078:begin
	ram_in<=32'd1008;
end
66079:begin
	ram_in<=32'd496;
end
66304:begin
	ram_in<=32'd32;
end
66305:begin
	ram_in<=32'd112;
end
66306:begin
	ram_in<=32'd496;
end
66307:begin
	ram_in<=32'd496;
end
66308:begin
	ram_in<=32'd1008;
end
66309:begin
	ram_in<=32'd1008;
end
66310:begin
	ram_in<=32'd496;
end
66311:begin
	ram_in<=32'd1008;
end
66312:begin
	ram_in<=32'd1008;
end
66313:begin
	ram_in<=32'd1008;
end
66314:begin
	ram_in<=32'd2032;
end
66315:begin
	ram_in<=32'd2032;
end
66316:begin
	ram_in<=32'd4064;
end
66317:begin
	ram_in<=32'd4080;
end
66318:begin
	ram_in<=32'd4080;
end
66319:begin
	ram_in<=32'd8176;
end
66320:begin
	ram_in<=32'd8176;
end
66321:begin
	ram_in<=32'd4064;
end
66322:begin
	ram_in<=32'd4064;
end
66323:begin
	ram_in<=32'd992;
end
66324:begin
	ram_in<=32'd496;
end
66325:begin
	ram_in<=32'd480;
end
66326:begin
	ram_in<=32'd480;
end
66327:begin
	ram_in<=32'd480;
end
66328:begin
	ram_in<=32'd480;
end
66329:begin
	ram_in<=32'd480;
end
66330:begin
	ram_in<=32'd992;
end
66331:begin
	ram_in<=32'd496;
end
66332:begin
	ram_in<=32'd496;
end
66333:begin
	ram_in<=32'd496;
end
66334:begin
	ram_in<=32'd496;
end
66335:begin
	ram_in<=32'd0;
end
66560:begin
	ram_in<=32'd192;
end
66561:begin
	ram_in<=32'd224;
end
66562:begin
	ram_in<=32'd1008;
end
66563:begin
	ram_in<=32'd496;
end
66564:begin
	ram_in<=32'd496;
end
66565:begin
	ram_in<=32'd496;
end
66566:begin
	ram_in<=32'd1008;
end
66567:begin
	ram_in<=32'd1008;
end
66568:begin
	ram_in<=32'd1008;
end
66569:begin
	ram_in<=32'd2016;
end
66570:begin
	ram_in<=32'd2016;
end
66571:begin
	ram_in<=32'd4032;
end
66572:begin
	ram_in<=32'd4064;
end
66573:begin
	ram_in<=32'd8160;
end
66574:begin
	ram_in<=32'd8160;
end
66575:begin
	ram_in<=32'd8128;
end
66576:begin
	ram_in<=32'd4032;
end
66577:begin
	ram_in<=32'd4032;
end
66578:begin
	ram_in<=32'd1984;
end
66579:begin
	ram_in<=32'd1984;
end
66580:begin
	ram_in<=32'd960;
end
66581:begin
	ram_in<=32'd960;
end
66582:begin
	ram_in<=32'd960;
end
66583:begin
	ram_in<=32'd960;
end
66584:begin
	ram_in<=32'd960;
end
66585:begin
	ram_in<=32'd992;
end
66586:begin
	ram_in<=32'd992;
end
66587:begin
	ram_in<=32'd992;
end
66588:begin
	ram_in<=32'd1008;
end
66589:begin
	ram_in<=32'd1008;
end
66590:begin
	ram_in<=32'd496;
end
66591:begin
	ram_in<=32'd32;
end
66816:begin
	ram_in<=32'd96;
end
66817:begin
	ram_in<=32'd240;
end
66818:begin
	ram_in<=32'd240;
end
66819:begin
	ram_in<=32'd240;
end
66820:begin
	ram_in<=32'd496;
end
66821:begin
	ram_in<=32'd496;
end
66822:begin
	ram_in<=32'd496;
end
66823:begin
	ram_in<=32'd1008;
end
66824:begin
	ram_in<=32'd1008;
end
66825:begin
	ram_in<=32'd2032;
end
66826:begin
	ram_in<=32'd2032;
end
66827:begin
	ram_in<=32'd2032;
end
66828:begin
	ram_in<=32'd4080;
end
66829:begin
	ram_in<=32'd4064;
end
66830:begin
	ram_in<=32'd8160;
end
66831:begin
	ram_in<=32'd8160;
end
66832:begin
	ram_in<=32'd4064;
end
66833:begin
	ram_in<=32'd992;
end
66834:begin
	ram_in<=32'd992;
end
66835:begin
	ram_in<=32'd992;
end
66836:begin
	ram_in<=32'd992;
end
66837:begin
	ram_in<=32'd992;
end
66838:begin
	ram_in<=32'd992;
end
66839:begin
	ram_in<=32'd496;
end
66840:begin
	ram_in<=32'd496;
end
66841:begin
	ram_in<=32'd496;
end
66842:begin
	ram_in<=32'd248;
end
66843:begin
	ram_in<=32'd508;
end
66844:begin
	ram_in<=32'd252;
end
66845:begin
	ram_in<=32'd252;
end
66846:begin
	ram_in<=32'd248;
end
66847:begin
	ram_in<=32'd112;
end
67072:begin
	ram_in<=32'd0;
end
67073:begin
	ram_in<=32'd960;
end
67074:begin
	ram_in<=32'd2016;
end
67075:begin
	ram_in<=32'd2016;
end
67076:begin
	ram_in<=32'd1008;
end
67077:begin
	ram_in<=32'd2032;
end
67078:begin
	ram_in<=32'd2032;
end
67079:begin
	ram_in<=32'd2032;
end
67080:begin
	ram_in<=32'd2032;
end
67081:begin
	ram_in<=32'd2032;
end
67082:begin
	ram_in<=32'd2032;
end
67083:begin
	ram_in<=32'd2032;
end
67084:begin
	ram_in<=32'd2032;
end
67085:begin
	ram_in<=32'd2016;
end
67086:begin
	ram_in<=32'd2032;
end
67087:begin
	ram_in<=32'd2016;
end
67088:begin
	ram_in<=32'd2016;
end
67089:begin
	ram_in<=32'd2016;
end
67090:begin
	ram_in<=32'd2032;
end
67091:begin
	ram_in<=32'd2032;
end
67092:begin
	ram_in<=32'd2016;
end
67093:begin
	ram_in<=32'd1984;
end
67094:begin
	ram_in<=32'd4064;
end
67095:begin
	ram_in<=32'd4064;
end
67096:begin
	ram_in<=32'd2016;
end
67097:begin
	ram_in<=32'd2016;
end
67098:begin
	ram_in<=32'd1984;
end
67099:begin
	ram_in<=32'd1984;
end
67100:begin
	ram_in<=32'd1984;
end
67101:begin
	ram_in<=32'd992;
end
67102:begin
	ram_in<=32'd224;
end
67103:begin
	ram_in<=32'd0;
end
67328:begin
	ram_in<=32'd0;
end
67329:begin
	ram_in<=32'd960;
end
67330:begin
	ram_in<=32'd992;
end
67331:begin
	ram_in<=32'd992;
end
67332:begin
	ram_in<=32'd1008;
end
67333:begin
	ram_in<=32'd1008;
end
67334:begin
	ram_in<=32'd1008;
end
67335:begin
	ram_in<=32'd1008;
end
67336:begin
	ram_in<=32'd1008;
end
67337:begin
	ram_in<=32'd1008;
end
67338:begin
	ram_in<=32'd992;
end
67339:begin
	ram_in<=32'd2016;
end
67340:begin
	ram_in<=32'd2016;
end
67341:begin
	ram_in<=32'd1008;
end
67342:begin
	ram_in<=32'd1008;
end
67343:begin
	ram_in<=32'd1008;
end
67344:begin
	ram_in<=32'd1008;
end
67345:begin
	ram_in<=32'd2032;
end
67346:begin
	ram_in<=32'd2016;
end
67347:begin
	ram_in<=32'd2016;
end
67348:begin
	ram_in<=32'd2016;
end
67349:begin
	ram_in<=32'd2016;
end
67350:begin
	ram_in<=32'd2016;
end
67351:begin
	ram_in<=32'd2016;
end
67352:begin
	ram_in<=32'd2016;
end
67353:begin
	ram_in<=32'd2016;
end
67354:begin
	ram_in<=32'd1008;
end
67355:begin
	ram_in<=32'd2032;
end
67356:begin
	ram_in<=32'd1008;
end
67357:begin
	ram_in<=32'd1008;
end
67358:begin
	ram_in<=32'd496;
end
67359:begin
	ram_in<=32'd0;
end
67584:begin
	ram_in<=32'd896;
end
67585:begin
	ram_in<=32'd1984;
end
67586:begin
	ram_in<=32'd2016;
end
67587:begin
	ram_in<=32'd2016;
end
67588:begin
	ram_in<=32'd2016;
end
67589:begin
	ram_in<=32'd2016;
end
67590:begin
	ram_in<=32'd2032;
end
67591:begin
	ram_in<=32'd4064;
end
67592:begin
	ram_in<=32'd4064;
end
67593:begin
	ram_in<=32'd1984;
end
67594:begin
	ram_in<=32'd4032;
end
67595:begin
	ram_in<=32'd4032;
end
67596:begin
	ram_in<=32'd1984;
end
67597:begin
	ram_in<=32'd1984;
end
67598:begin
	ram_in<=32'd4032;
end
67599:begin
	ram_in<=32'd4064;
end
67600:begin
	ram_in<=32'd4064;
end
67601:begin
	ram_in<=32'd4064;
end
67602:begin
	ram_in<=32'd2016;
end
67603:begin
	ram_in<=32'd4032;
end
67604:begin
	ram_in<=32'd1984;
end
67605:begin
	ram_in<=32'd2016;
end
67606:begin
	ram_in<=32'd4064;
end
67607:begin
	ram_in<=32'd4064;
end
67608:begin
	ram_in<=32'd2016;
end
67609:begin
	ram_in<=32'd2016;
end
67610:begin
	ram_in<=32'd2016;
end
67611:begin
	ram_in<=32'd2032;
end
67612:begin
	ram_in<=32'd2032;
end
67613:begin
	ram_in<=32'd2032;
end
67614:begin
	ram_in<=32'd192;
end
67615:begin
	ram_in<=32'd128;
end
67840:begin
	ram_in<=32'd16;
end
67841:begin
	ram_in<=32'd56;
end
67842:begin
	ram_in<=32'd56;
end
67843:begin
	ram_in<=32'd56;
end
67844:begin
	ram_in<=32'd120;
end
67845:begin
	ram_in<=32'd120;
end
67846:begin
	ram_in<=32'd120;
end
67847:begin
	ram_in<=32'd248;
end
67848:begin
	ram_in<=32'd504;
end
67849:begin
	ram_in<=32'd1008;
end
67850:begin
	ram_in<=32'd2032;
end
67851:begin
	ram_in<=32'd2032;
end
67852:begin
	ram_in<=32'd4080;
end
67853:begin
	ram_in<=32'd4080;
end
67854:begin
	ram_in<=32'd8176;
end
67855:begin
	ram_in<=32'd7920;
end
67856:begin
	ram_in<=32'd7408;
end
67857:begin
	ram_in<=32'd3312;
end
67858:begin
	ram_in<=32'd1136;
end
67859:begin
	ram_in<=32'd112;
end
67860:begin
	ram_in<=32'd240;
end
67861:begin
	ram_in<=32'd240;
end
67862:begin
	ram_in<=32'd240;
end
67863:begin
	ram_in<=32'd112;
end
67864:begin
	ram_in<=32'd112;
end
67865:begin
	ram_in<=32'd112;
end
67866:begin
	ram_in<=32'd56;
end
67867:begin
	ram_in<=32'd112;
end
67868:begin
	ram_in<=32'd112;
end
67869:begin
	ram_in<=32'd48;
end
67870:begin
	ram_in<=32'd48;
end
67871:begin
	ram_in<=32'd48;
end
131072:begin
	ram_in<=32'd1792;
end
131073:begin
	ram_in<=32'd3968;
end
131074:begin
	ram_in<=32'd8064;
end
131075:begin
	ram_in<=32'd4032;
end
131076:begin
	ram_in<=32'd4032;
end
131077:begin
	ram_in<=32'd4032;
end
131078:begin
	ram_in<=32'd3552;
end
131079:begin
	ram_in<=32'd3296;
end
131080:begin
	ram_in<=32'd3296;
end
131081:begin
	ram_in<=32'd2272;
end
131082:begin
	ram_in<=32'd2272;
end
131083:begin
	ram_in<=32'd192;
end
131084:begin
	ram_in<=32'd224;
end
131085:begin
	ram_in<=32'd224;
end
131086:begin
	ram_in<=32'd224;
end
131087:begin
	ram_in<=32'd224;
end
131088:begin
	ram_in<=32'd224;
end
131089:begin
	ram_in<=32'd448;
end
131090:begin
	ram_in<=32'd448;
end
131091:begin
	ram_in<=32'd448;
end
131092:begin
	ram_in<=32'd896;
end
131093:begin
	ram_in<=32'd448;
end
131094:begin
	ram_in<=32'd960;
end
131095:begin
	ram_in<=32'd1920;
end
131096:begin
	ram_in<=32'd1920;
end
131097:begin
	ram_in<=32'd4092;
end
131098:begin
	ram_in<=32'd4092;
end
131099:begin
	ram_in<=32'd8188;
end
131100:begin
	ram_in<=32'd8188;
end
131101:begin
	ram_in<=32'd8188;
end
131102:begin
	ram_in<=32'd4092;
end
131103:begin
	ram_in<=32'd4032;
end
131328:begin
	ram_in<=32'd768;
end
131329:begin
	ram_in<=32'd896;
end
131330:begin
	ram_in<=32'd1920;
end
131331:begin
	ram_in<=32'd1984;
end
131332:begin
	ram_in<=32'd4032;
end
131333:begin
	ram_in<=32'd1984;
end
131334:begin
	ram_in<=32'd3776;
end
131335:begin
	ram_in<=32'd3776;
end
131336:begin
	ram_in<=32'd3680;
end
131337:begin
	ram_in<=32'd3136;
end
131338:begin
	ram_in<=32'd3136;
end
131339:begin
	ram_in<=32'd3168;
end
131340:begin
	ram_in<=32'd3168;
end
131341:begin
	ram_in<=32'd3168;
end
131342:begin
	ram_in<=32'd3264;
end
131343:begin
	ram_in<=32'd1120;
end
131344:begin
	ram_in<=32'd64;
end
131345:begin
	ram_in<=32'd192;
end
131346:begin
	ram_in<=32'd224;
end
131347:begin
	ram_in<=32'd192;
end
131348:begin
	ram_in<=32'd448;
end
131349:begin
	ram_in<=32'd448;
end
131350:begin
	ram_in<=32'd192;
end
131351:begin
	ram_in<=32'd448;
end
131352:begin
	ram_in<=32'd1016;
end
131353:begin
	ram_in<=32'd1022;
end
131354:begin
	ram_in<=32'd2046;
end
131355:begin
	ram_in<=32'd2046;
end
131356:begin
	ram_in<=32'd2046;
end
131357:begin
	ram_in<=32'd2046;
end
131358:begin
	ram_in<=32'd768;
end
131359:begin
	ram_in<=32'd0;
end
131584:begin
	ram_in<=32'd512;
end
131585:begin
	ram_in<=32'd896;
end
131586:begin
	ram_in<=32'd1984;
end
131587:begin
	ram_in<=32'd4032;
end
131588:begin
	ram_in<=32'd4032;
end
131589:begin
	ram_in<=32'd4064;
end
131590:begin
	ram_in<=32'd8160;
end
131591:begin
	ram_in<=32'd7392;
end
131592:begin
	ram_in<=32'd2144;
end
131593:begin
	ram_in<=32'd2144;
end
131594:begin
	ram_in<=32'd96;
end
131595:begin
	ram_in<=32'd96;
end
131596:begin
	ram_in<=32'd96;
end
131597:begin
	ram_in<=32'd96;
end
131598:begin
	ram_in<=32'd96;
end
131599:begin
	ram_in<=32'd96;
end
131600:begin
	ram_in<=32'd96;
end
131601:begin
	ram_in<=32'd224;
end
131602:begin
	ram_in<=32'd224;
end
131603:begin
	ram_in<=32'd192;
end
131604:begin
	ram_in<=32'd448;
end
131605:begin
	ram_in<=32'd448;
end
131606:begin
	ram_in<=32'd896;
end
131607:begin
	ram_in<=32'd896;
end
131608:begin
	ram_in<=32'd896;
end
131609:begin
	ram_in<=32'd2040;
end
131610:begin
	ram_in<=32'd2040;
end
131611:begin
	ram_in<=32'd4088;
end
131612:begin
	ram_in<=32'd2040;
end
131613:begin
	ram_in<=32'd2040;
end
131614:begin
	ram_in<=32'd4064;
end
131615:begin
	ram_in<=32'd0;
end
131840:begin
	ram_in<=32'd256;
end
131841:begin
	ram_in<=32'd384;
end
131842:begin
	ram_in<=32'd1984;
end
131843:begin
	ram_in<=32'd4032;
end
131844:begin
	ram_in<=32'd4032;
end
131845:begin
	ram_in<=32'd4032;
end
131846:begin
	ram_in<=32'd8160;
end
131847:begin
	ram_in<=32'd7392;
end
131848:begin
	ram_in<=32'd7264;
end
131849:begin
	ram_in<=32'd6240;
end
131850:begin
	ram_in<=32'd6240;
end
131851:begin
	ram_in<=32'd6240;
end
131852:begin
	ram_in<=32'd64;
end
131853:begin
	ram_in<=32'd96;
end
131854:begin
	ram_in<=32'd96;
end
131855:begin
	ram_in<=32'd96;
end
131856:begin
	ram_in<=32'd96;
end
131857:begin
	ram_in<=32'd192;
end
131858:begin
	ram_in<=32'd192;
end
131859:begin
	ram_in<=32'd192;
end
131860:begin
	ram_in<=32'd192;
end
131861:begin
	ram_in<=32'd192;
end
131862:begin
	ram_in<=32'd448;
end
131863:begin
	ram_in<=32'd384;
end
131864:begin
	ram_in<=32'd992;
end
131865:begin
	ram_in<=32'd1016;
end
131866:begin
	ram_in<=32'd4092;
end
131867:begin
	ram_in<=32'd2044;
end
131868:begin
	ram_in<=32'd2044;
end
131869:begin
	ram_in<=32'd2044;
end
131870:begin
	ram_in<=32'd4036;
end
131871:begin
	ram_in<=32'd512;
end
132096:begin
	ram_in<=32'd896;
end
132097:begin
	ram_in<=32'd896;
end
132098:begin
	ram_in<=32'd4032;
end
132099:begin
	ram_in<=32'd4032;
end
132100:begin
	ram_in<=32'd4032;
end
132101:begin
	ram_in<=32'd8160;
end
132102:begin
	ram_in<=32'd3696;
end
132103:begin
	ram_in<=32'd3168;
end
132104:begin
	ram_in<=32'd2144;
end
132105:begin
	ram_in<=32'd2144;
end
132106:begin
	ram_in<=32'd96;
end
132107:begin
	ram_in<=32'd96;
end
132108:begin
	ram_in<=32'd96;
end
132109:begin
	ram_in<=32'd96;
end
132110:begin
	ram_in<=32'd96;
end
132111:begin
	ram_in<=32'd224;
end
132112:begin
	ram_in<=32'd192;
end
132113:begin
	ram_in<=32'd192;
end
132114:begin
	ram_in<=32'd192;
end
132115:begin
	ram_in<=32'd448;
end
132116:begin
	ram_in<=32'd192;
end
132117:begin
	ram_in<=32'd448;
end
132118:begin
	ram_in<=32'd384;
end
132119:begin
	ram_in<=32'd896;
end
132120:begin
	ram_in<=32'd896;
end
132121:begin
	ram_in<=32'd1848;
end
132122:begin
	ram_in<=32'd4088;
end
132123:begin
	ram_in<=32'd2044;
end
132124:begin
	ram_in<=32'd2044;
end
132125:begin
	ram_in<=32'd4092;
end
132126:begin
	ram_in<=32'd4092;
end
132127:begin
	ram_in<=32'd8;
end
132352:begin
	ram_in<=32'd1536;
end
132353:begin
	ram_in<=32'd1792;
end
132354:begin
	ram_in<=32'd3840;
end
132355:begin
	ram_in<=32'd3968;
end
132356:begin
	ram_in<=32'd8128;
end
132357:begin
	ram_in<=32'd8128;
end
132358:begin
	ram_in<=32'd8128;
end
132359:begin
	ram_in<=32'd7616;
end
132360:begin
	ram_in<=32'd7360;
end
132361:begin
	ram_in<=32'd7360;
end
132362:begin
	ram_in<=32'd2240;
end
132363:begin
	ram_in<=32'd224;
end
132364:begin
	ram_in<=32'd224;
end
132365:begin
	ram_in<=32'd192;
end
132366:begin
	ram_in<=32'd224;
end
132367:begin
	ram_in<=32'd224;
end
132368:begin
	ram_in<=32'd192;
end
132369:begin
	ram_in<=32'd448;
end
132370:begin
	ram_in<=32'd448;
end
132371:begin
	ram_in<=32'd448;
end
132372:begin
	ram_in<=32'd448;
end
132373:begin
	ram_in<=32'd448;
end
132374:begin
	ram_in<=32'd896;
end
132375:begin
	ram_in<=32'd1920;
end
132376:begin
	ram_in<=32'd3984;
end
132377:begin
	ram_in<=32'd2044;
end
132378:begin
	ram_in<=32'd4092;
end
132379:begin
	ram_in<=32'd4092;
end
132380:begin
	ram_in<=32'd4092;
end
132381:begin
	ram_in<=32'd4092;
end
132382:begin
	ram_in<=32'd2046;
end
132383:begin
	ram_in<=32'd46;
end
132608:begin
	ram_in<=32'd512;
end
132609:begin
	ram_in<=32'd1920;
end
132610:begin
	ram_in<=32'd4032;
end
132611:begin
	ram_in<=32'd3008;
end
132612:begin
	ram_in<=32'd3008;
end
132613:begin
	ram_in<=32'd4032;
end
132614:begin
	ram_in<=32'd8160;
end
132615:begin
	ram_in<=32'd7776;
end
132616:begin
	ram_in<=32'd2144;
end
132617:begin
	ram_in<=32'd96;
end
132618:begin
	ram_in<=32'd112;
end
132619:begin
	ram_in<=32'd96;
end
132620:begin
	ram_in<=32'd96;
end
132621:begin
	ram_in<=32'd96;
end
132622:begin
	ram_in<=32'd96;
end
132623:begin
	ram_in<=32'd96;
end
132624:begin
	ram_in<=32'd96;
end
132625:begin
	ram_in<=32'd96;
end
132626:begin
	ram_in<=32'd96;
end
132627:begin
	ram_in<=32'd192;
end
132628:begin
	ram_in<=32'd192;
end
132629:begin
	ram_in<=32'd448;
end
132630:begin
	ram_in<=32'd448;
end
132631:begin
	ram_in<=32'd384;
end
132632:begin
	ram_in<=32'd896;
end
132633:begin
	ram_in<=32'd1936;
end
132634:begin
	ram_in<=32'd2040;
end
132635:begin
	ram_in<=32'd2040;
end
132636:begin
	ram_in<=32'd2040;
end
132637:begin
	ram_in<=32'd4088;
end
132638:begin
	ram_in<=32'd4088;
end
132639:begin
	ram_in<=32'd504;
end
132864:begin
	ram_in<=32'd896;
end
132865:begin
	ram_in<=32'd1920;
end
132866:begin
	ram_in<=32'd3968;
end
132867:begin
	ram_in<=32'd1984;
end
132868:begin
	ram_in<=32'd4032;
end
132869:begin
	ram_in<=32'd4032;
end
132870:begin
	ram_in<=32'd4032;
end
132871:begin
	ram_in<=32'd4064;
end
132872:begin
	ram_in<=32'd3808;
end
132873:begin
	ram_in<=32'd1248;
end
132874:begin
	ram_in<=32'd1248;
end
132875:begin
	ram_in<=32'd96;
end
132876:begin
	ram_in<=32'd96;
end
132877:begin
	ram_in<=32'd224;
end
132878:begin
	ram_in<=32'd224;
end
132879:begin
	ram_in<=32'd112;
end
132880:begin
	ram_in<=32'd224;
end
132881:begin
	ram_in<=32'd224;
end
132882:begin
	ram_in<=32'd240;
end
132883:begin
	ram_in<=32'd240;
end
132884:begin
	ram_in<=32'd240;
end
132885:begin
	ram_in<=32'd504;
end
132886:begin
	ram_in<=32'd508;
end
132887:begin
	ram_in<=32'd1020;
end
132888:begin
	ram_in<=32'd1020;
end
132889:begin
	ram_in<=32'd2046;
end
132890:begin
	ram_in<=32'd2046;
end
132891:begin
	ram_in<=32'd1990;
end
132892:begin
	ram_in<=32'd3974;
end
132893:begin
	ram_in<=32'd3846;
end
132894:begin
	ram_in<=32'd1794;
end
132895:begin
	ram_in<=32'd1792;
end
133120:begin
	ram_in<=32'd448;
end
133121:begin
	ram_in<=32'd2016;
end
133122:begin
	ram_in<=32'd2016;
end
133123:begin
	ram_in<=32'd4080;
end
133124:begin
	ram_in<=32'd4080;
end
133125:begin
	ram_in<=32'd3704;
end
133126:begin
	ram_in<=32'd3120;
end
133127:begin
	ram_in<=32'd2104;
end
133128:begin
	ram_in<=32'd56;
end
133129:begin
	ram_in<=32'd56;
end
133130:begin
	ram_in<=32'd112;
end
133131:begin
	ram_in<=32'd224;
end
133132:begin
	ram_in<=32'd224;
end
133133:begin
	ram_in<=32'd224;
end
133134:begin
	ram_in<=32'd448;
end
133135:begin
	ram_in<=32'd448;
end
133136:begin
	ram_in<=32'd896;
end
133137:begin
	ram_in<=32'd256;
end
133138:begin
	ram_in<=32'd1792;
end
133139:begin
	ram_in<=32'd1536;
end
133140:begin
	ram_in<=32'd3584;
end
133141:begin
	ram_in<=32'd1536;
end
133142:begin
	ram_in<=32'd3072;
end
133143:begin
	ram_in<=32'd7168;
end
133144:begin
	ram_in<=32'd6144;
end
133145:begin
	ram_in<=32'd7616;
end
133146:begin
	ram_in<=32'd8176;
end
133147:begin
	ram_in<=32'd8184;
end
133148:begin
	ram_in<=32'd4088;
end
133149:begin
	ram_in<=32'd2040;
end
133150:begin
	ram_in<=32'd24;
end
133151:begin
	ram_in<=32'd8;
end
133376:begin
	ram_in<=32'd1536;
end
133377:begin
	ram_in<=32'd3840;
end
133378:begin
	ram_in<=32'd3840;
end
133379:begin
	ram_in<=32'd8064;
end
133380:begin
	ram_in<=32'd8064;
end
133381:begin
	ram_in<=32'd8128;
end
133382:begin
	ram_in<=32'd8128;
end
133383:begin
	ram_in<=32'd6336;
end
133384:begin
	ram_in<=32'd6336;
end
133385:begin
	ram_in<=32'd6336;
end
133386:begin
	ram_in<=32'd4288;
end
133387:begin
	ram_in<=32'd192;
end
133388:begin
	ram_in<=32'd192;
end
133389:begin
	ram_in<=32'd192;
end
133390:begin
	ram_in<=32'd192;
end
133391:begin
	ram_in<=32'd448;
end
133392:begin
	ram_in<=32'd448;
end
133393:begin
	ram_in<=32'd384;
end
133394:begin
	ram_in<=32'd896;
end
133395:begin
	ram_in<=32'd896;
end
133396:begin
	ram_in<=32'd768;
end
133397:begin
	ram_in<=32'd896;
end
133398:begin
	ram_in<=32'd768;
end
133399:begin
	ram_in<=32'd1792;
end
133400:begin
	ram_in<=32'd1584;
end
133401:begin
	ram_in<=32'd2040;
end
133402:begin
	ram_in<=32'd4092;
end
133403:begin
	ram_in<=32'd4092;
end
133404:begin
	ram_in<=32'd4092;
end
133405:begin
	ram_in<=32'd4088;
end
133406:begin
	ram_in<=32'd2032;
end
133407:begin
	ram_in<=32'd1536;
end
196608:begin
	ram_in<=32'd448;
end
196609:begin
	ram_in<=32'd1984;
end
196610:begin
	ram_in<=32'd4064;
end
196611:begin
	ram_in<=32'd2032;
end
196612:begin
	ram_in<=32'd4080;
end
196613:begin
	ram_in<=32'd4080;
end
196614:begin
	ram_in<=32'd3632;
end
196615:begin
	ram_in<=32'd3120;
end
196616:begin
	ram_in<=32'd112;
end
196617:begin
	ram_in<=32'd112;
end
196618:begin
	ram_in<=32'd240;
end
196619:begin
	ram_in<=32'd224;
end
196620:begin
	ram_in<=32'd480;
end
196621:begin
	ram_in<=32'd960;
end
196622:begin
	ram_in<=32'd992;
end
196623:begin
	ram_in<=32'd992;
end
196624:begin
	ram_in<=32'd992;
end
196625:begin
	ram_in<=32'd1008;
end
196626:begin
	ram_in<=32'd1008;
end
196627:begin
	ram_in<=32'd56;
end
196628:begin
	ram_in<=32'd24;
end
196629:begin
	ram_in<=32'd24;
end
196630:begin
	ram_in<=32'd24;
end
196631:begin
	ram_in<=32'd28;
end
196632:begin
	ram_in<=32'd3612;
end
196633:begin
	ram_in<=32'd1564;
end
196634:begin
	ram_in<=32'd1596;
end
196635:begin
	ram_in<=32'd4088;
end
196636:begin
	ram_in<=32'd2040;
end
196637:begin
	ram_in<=32'd4080;
end
196638:begin
	ram_in<=32'd2032;
end
196639:begin
	ram_in<=32'd992;
end
196864:begin
	ram_in<=32'd448;
end
196865:begin
	ram_in<=32'd960;
end
196866:begin
	ram_in<=32'd4032;
end
196867:begin
	ram_in<=32'd2016;
end
196868:begin
	ram_in<=32'd1904;
end
196869:begin
	ram_in<=32'd1648;
end
196870:begin
	ram_in<=32'd1072;
end
196871:begin
	ram_in<=32'd48;
end
196872:begin
	ram_in<=32'd48;
end
196873:begin
	ram_in<=32'd112;
end
196874:begin
	ram_in<=32'd96;
end
196875:begin
	ram_in<=32'd224;
end
196876:begin
	ram_in<=32'd992;
end
196877:begin
	ram_in<=32'd992;
end
196878:begin
	ram_in<=32'd992;
end
196879:begin
	ram_in<=32'd992;
end
196880:begin
	ram_in<=32'd992;
end
196881:begin
	ram_in<=32'd1008;
end
196882:begin
	ram_in<=32'd240;
end
196883:begin
	ram_in<=32'd48;
end
196884:begin
	ram_in<=32'd24;
end
196885:begin
	ram_in<=32'd28;
end
196886:begin
	ram_in<=32'd12;
end
196887:begin
	ram_in<=32'd12;
end
196888:begin
	ram_in<=32'd1052;
end
196889:begin
	ram_in<=32'd3100;
end
196890:begin
	ram_in<=32'd3640;
end
196891:begin
	ram_in<=32'd3704;
end
196892:begin
	ram_in<=32'd4088;
end
196893:begin
	ram_in<=32'd4080;
end
196894:begin
	ram_in<=32'd2032;
end
196895:begin
	ram_in<=32'd960;
end
197120:begin
	ram_in<=32'd0;
end
197121:begin
	ram_in<=32'd960;
end
197122:begin
	ram_in<=32'd1984;
end
197123:begin
	ram_in<=32'd4064;
end
197124:begin
	ram_in<=32'd4064;
end
197125:begin
	ram_in<=32'd7264;
end
197126:begin
	ram_in<=32'd7216;
end
197127:begin
	ram_in<=32'd6192;
end
197128:begin
	ram_in<=32'd6192;
end
197129:begin
	ram_in<=32'd6240;
end
197130:begin
	ram_in<=32'd4192;
end
197131:begin
	ram_in<=32'd224;
end
197132:begin
	ram_in<=32'd224;
end
197133:begin
	ram_in<=32'd192;
end
197134:begin
	ram_in<=32'd448;
end
197135:begin
	ram_in<=32'd2016;
end
197136:begin
	ram_in<=32'd2016;
end
197137:begin
	ram_in<=32'd2032;
end
197138:begin
	ram_in<=32'd2032;
end
197139:begin
	ram_in<=32'd56;
end
197140:begin
	ram_in<=32'd28;
end
197141:begin
	ram_in<=32'd12;
end
197142:begin
	ram_in<=32'd12;
end
197143:begin
	ram_in<=32'd12;
end
197144:begin
	ram_in<=32'd12;
end
197145:begin
	ram_in<=32'd3100;
end
197146:begin
	ram_in<=32'd3640;
end
197147:begin
	ram_in<=32'd2040;
end
197148:begin
	ram_in<=32'd2040;
end
197149:begin
	ram_in<=32'd2032;
end
197150:begin
	ram_in<=32'd992;
end
197151:begin
	ram_in<=32'd128;
end
197376:begin
	ram_in<=32'd192;
end
197377:begin
	ram_in<=32'd992;
end
197378:begin
	ram_in<=32'd4080;
end
197379:begin
	ram_in<=32'd4080;
end
197380:begin
	ram_in<=32'd8184;
end
197381:begin
	ram_in<=32'd7728;
end
197382:begin
	ram_in<=32'd7216;
end
197383:begin
	ram_in<=32'd6256;
end
197384:begin
	ram_in<=32'd6240;
end
197385:begin
	ram_in<=32'd224;
end
197386:begin
	ram_in<=32'd992;
end
197387:begin
	ram_in<=32'd960;
end
197388:begin
	ram_in<=32'd1984;
end
197389:begin
	ram_in<=32'd4032;
end
197390:begin
	ram_in<=32'd4064;
end
197391:begin
	ram_in<=32'd4064;
end
197392:begin
	ram_in<=32'd4080;
end
197393:begin
	ram_in<=32'd3184;
end
197394:begin
	ram_in<=32'd112;
end
197395:begin
	ram_in<=32'd56;
end
197396:begin
	ram_in<=32'd56;
end
197397:begin
	ram_in<=32'd24;
end
197398:begin
	ram_in<=32'd24;
end
197399:begin
	ram_in<=32'd24;
end
197400:begin
	ram_in<=32'd1592;
end
197401:begin
	ram_in<=32'd3632;
end
197402:begin
	ram_in<=32'd3824;
end
197403:begin
	ram_in<=32'd4080;
end
197404:begin
	ram_in<=32'd4064;
end
197405:begin
	ram_in<=32'd4064;
end
197406:begin
	ram_in<=32'd2016;
end
197407:begin
	ram_in<=32'd128;
end
197632:begin
	ram_in<=32'd768;
end
197633:begin
	ram_in<=32'd1920;
end
197634:begin
	ram_in<=32'd8064;
end
197635:begin
	ram_in<=32'd4032;
end
197636:begin
	ram_in<=32'd8128;
end
197637:begin
	ram_in<=32'd8128;
end
197638:begin
	ram_in<=32'd3264;
end
197639:begin
	ram_in<=32'd2240;
end
197640:begin
	ram_in<=32'd192;
end
197641:begin
	ram_in<=32'd448;
end
197642:begin
	ram_in<=32'd448;
end
197643:begin
	ram_in<=32'd960;
end
197644:begin
	ram_in<=32'd1920;
end
197645:begin
	ram_in<=32'd1920;
end
197646:begin
	ram_in<=32'd1792;
end
197647:begin
	ram_in<=32'd1792;
end
197648:begin
	ram_in<=32'd2032;
end
197649:begin
	ram_in<=32'd2032;
end
197650:begin
	ram_in<=32'd2040;
end
197651:begin
	ram_in<=32'd1016;
end
197652:begin
	ram_in<=32'd120;
end
197653:begin
	ram_in<=32'd24;
end
197654:begin
	ram_in<=32'd24;
end
197655:begin
	ram_in<=32'd24;
end
197656:begin
	ram_in<=32'd24;
end
197657:begin
	ram_in<=32'd120;
end
197658:begin
	ram_in<=32'd504;
end
197659:begin
	ram_in<=32'd2032;
end
197660:begin
	ram_in<=32'd8176;
end
197661:begin
	ram_in<=32'd8128;
end
197662:begin
	ram_in<=32'd4032;
end
197663:begin
	ram_in<=32'd0;
end
197888:begin
	ram_in<=32'd448;
end
197889:begin
	ram_in<=32'd2032;
end
197890:begin
	ram_in<=32'd4080;
end
197891:begin
	ram_in<=32'd4088;
end
197892:begin
	ram_in<=32'd4088;
end
197893:begin
	ram_in<=32'd3640;
end
197894:begin
	ram_in<=32'd2104;
end
197895:begin
	ram_in<=32'd56;
end
197896:begin
	ram_in<=32'd48;
end
197897:begin
	ram_in<=32'd48;
end
197898:begin
	ram_in<=32'd240;
end
197899:begin
	ram_in<=32'd224;
end
197900:begin
	ram_in<=32'd224;
end
197901:begin
	ram_in<=32'd448;
end
197902:begin
	ram_in<=32'd448;
end
197903:begin
	ram_in<=32'd448;
end
197904:begin
	ram_in<=32'd480;
end
197905:begin
	ram_in<=32'd496;
end
197906:begin
	ram_in<=32'd248;
end
197907:begin
	ram_in<=32'd248;
end
197908:begin
	ram_in<=32'd120;
end
197909:begin
	ram_in<=32'd56;
end
197910:begin
	ram_in<=32'd24;
end
197911:begin
	ram_in<=32'd24;
end
197912:begin
	ram_in<=32'd24;
end
197913:begin
	ram_in<=32'd2104;
end
197914:begin
	ram_in<=32'd6264;
end
197915:begin
	ram_in<=32'd8184;
end
197916:begin
	ram_in<=32'd8176;
end
197917:begin
	ram_in<=32'd4080;
end
197918:begin
	ram_in<=32'd4064;
end
197919:begin
	ram_in<=32'd640;
end
198144:begin
	ram_in<=32'd128;
end
198145:begin
	ram_in<=32'd992;
end
198146:begin
	ram_in<=32'd4080;
end
198147:begin
	ram_in<=32'd4064;
end
198148:begin
	ram_in<=32'd8176;
end
198149:begin
	ram_in<=32'd8048;
end
198150:begin
	ram_in<=32'd7216;
end
198151:begin
	ram_in<=32'd2096;
end
198152:begin
	ram_in<=32'd2096;
end
198153:begin
	ram_in<=32'd48;
end
198154:begin
	ram_in<=32'd112;
end
198155:begin
	ram_in<=32'd96;
end
198156:begin
	ram_in<=32'd224;
end
198157:begin
	ram_in<=32'd224;
end
198158:begin
	ram_in<=32'd480;
end
198159:begin
	ram_in<=32'd448;
end
198160:begin
	ram_in<=32'd480;
end
198161:begin
	ram_in<=32'd480;
end
198162:begin
	ram_in<=32'd224;
end
198163:begin
	ram_in<=32'd240;
end
198164:begin
	ram_in<=32'd120;
end
198165:begin
	ram_in<=32'd56;
end
198166:begin
	ram_in<=32'd24;
end
198167:begin
	ram_in<=32'd24;
end
198168:begin
	ram_in<=32'd24;
end
198169:begin
	ram_in<=32'd2072;
end
198170:begin
	ram_in<=32'd2168;
end
198171:begin
	ram_in<=32'd4088;
end
198172:begin
	ram_in<=32'd4088;
end
198173:begin
	ram_in<=32'd4080;
end
198174:begin
	ram_in<=32'd4064;
end
198175:begin
	ram_in<=32'd384;
end
198400:begin
	ram_in<=32'd832;
end
198401:begin
	ram_in<=32'd2016;
end
198402:begin
	ram_in<=32'd4064;
end
198403:begin
	ram_in<=32'd8160;
end
198404:begin
	ram_in<=32'd8160;
end
198405:begin
	ram_in<=32'd8160;
end
198406:begin
	ram_in<=32'd4064;
end
198407:begin
	ram_in<=32'd224;
end
198408:begin
	ram_in<=32'd224;
end
198409:begin
	ram_in<=32'd224;
end
198410:begin
	ram_in<=32'd224;
end
198411:begin
	ram_in<=32'd448;
end
198412:begin
	ram_in<=32'd448;
end
198413:begin
	ram_in<=32'd448;
end
198414:begin
	ram_in<=32'd448;
end
198415:begin
	ram_in<=32'd480;
end
198416:begin
	ram_in<=32'd496;
end
198417:begin
	ram_in<=32'd240;
end
198418:begin
	ram_in<=32'd248;
end
198419:begin
	ram_in<=32'd120;
end
198420:begin
	ram_in<=32'd56;
end
198421:begin
	ram_in<=32'd24;
end
198422:begin
	ram_in<=32'd24;
end
198423:begin
	ram_in<=32'd24;
end
198424:begin
	ram_in<=32'd24;
end
198425:begin
	ram_in<=32'd24;
end
198426:begin
	ram_in<=32'd3192;
end
198427:begin
	ram_in<=32'd4088;
end
198428:begin
	ram_in<=32'd4080;
end
198429:begin
	ram_in<=32'd4080;
end
198430:begin
	ram_in<=32'd4064;
end
198431:begin
	ram_in<=32'd896;
end
198656:begin
	ram_in<=32'd256;
end
198657:begin
	ram_in<=32'd896;
end
198658:begin
	ram_in<=32'd1984;
end
198659:begin
	ram_in<=32'd1984;
end
198660:begin
	ram_in<=32'd2016;
end
198661:begin
	ram_in<=32'd4064;
end
198662:begin
	ram_in<=32'd3296;
end
198663:begin
	ram_in<=32'd2144;
end
198664:begin
	ram_in<=32'd2144;
end
198665:begin
	ram_in<=32'd2144;
end
198666:begin
	ram_in<=32'd96;
end
198667:begin
	ram_in<=32'd96;
end
198668:begin
	ram_in<=32'd96;
end
198669:begin
	ram_in<=32'd192;
end
198670:begin
	ram_in<=32'd1984;
end
198671:begin
	ram_in<=32'd2016;
end
198672:begin
	ram_in<=32'd2016;
end
198673:begin
	ram_in<=32'd2016;
end
198674:begin
	ram_in<=32'd2032;
end
198675:begin
	ram_in<=32'd1904;
end
198676:begin
	ram_in<=32'd48;
end
198677:begin
	ram_in<=32'd48;
end
198678:begin
	ram_in<=32'd16;
end
198679:begin
	ram_in<=32'd24;
end
198680:begin
	ram_in<=32'd24;
end
198681:begin
	ram_in<=32'd536;
end
198682:begin
	ram_in<=32'd792;
end
198683:begin
	ram_in<=32'd2032;
end
198684:begin
	ram_in<=32'd2032;
end
198685:begin
	ram_in<=32'd2032;
end
198686:begin
	ram_in<=32'd992;
end
198687:begin
	ram_in<=32'd0;
end
198912:begin
	ram_in<=32'd64;
end
198913:begin
	ram_in<=32'd224;
end
198914:begin
	ram_in<=32'd1008;
end
198915:begin
	ram_in<=32'd2032;
end
198916:begin
	ram_in<=32'd2032;
end
198917:begin
	ram_in<=32'd2032;
end
198918:begin
	ram_in<=32'd4080;
end
198919:begin
	ram_in<=32'd1968;
end
198920:begin
	ram_in<=32'd3184;
end
198921:begin
	ram_in<=32'd3184;
end
198922:begin
	ram_in<=32'd1248;
end
198923:begin
	ram_in<=32'd224;
end
198924:begin
	ram_in<=32'd224;
end
198925:begin
	ram_in<=32'd224;
end
198926:begin
	ram_in<=32'd480;
end
198927:begin
	ram_in<=32'd480;
end
198928:begin
	ram_in<=32'd496;
end
198929:begin
	ram_in<=32'd240;
end
198930:begin
	ram_in<=32'd120;
end
198931:begin
	ram_in<=32'd112;
end
198932:begin
	ram_in<=32'd56;
end
198933:begin
	ram_in<=32'd24;
end
198934:begin
	ram_in<=32'd24;
end
198935:begin
	ram_in<=32'd24;
end
198936:begin
	ram_in<=32'd824;
end
198937:begin
	ram_in<=32'd624;
end
198938:begin
	ram_in<=32'd1008;
end
198939:begin
	ram_in<=32'd1008;
end
198940:begin
	ram_in<=32'd992;
end
198941:begin
	ram_in<=32'd960;
end
198942:begin
	ram_in<=32'd896;
end
198943:begin
	ram_in<=32'd768;
end
262144:begin
	ram_in<=32'd96;
end
262145:begin
	ram_in<=32'd112;
end
262146:begin
	ram_in<=32'd240;
end
262147:begin
	ram_in<=32'd240;
end
262148:begin
	ram_in<=32'd496;
end
262149:begin
	ram_in<=32'd1008;
end
262150:begin
	ram_in<=32'd2032;
end
262151:begin
	ram_in<=32'd1968;
end
262152:begin
	ram_in<=32'd1840;
end
262153:begin
	ram_in<=32'd3952;
end
262154:begin
	ram_in<=32'd3696;
end
262155:begin
	ram_in<=32'd7280;
end
262156:begin
	ram_in<=32'd7288;
end
262157:begin
	ram_in<=32'd7416;
end
262158:begin
	ram_in<=32'd8188;
end
262159:begin
	ram_in<=32'd8188;
end
262160:begin
	ram_in<=32'd8188;
end
262161:begin
	ram_in<=32'd8184;
end
262162:begin
	ram_in<=32'd8176;
end
262163:begin
	ram_in<=32'd3696;
end
262164:begin
	ram_in<=32'd96;
end
262165:begin
	ram_in<=32'd96;
end
262166:begin
	ram_in<=32'd96;
end
262167:begin
	ram_in<=32'd96;
end
262168:begin
	ram_in<=32'd96;
end
262169:begin
	ram_in<=32'd96;
end
262170:begin
	ram_in<=32'd96;
end
262171:begin
	ram_in<=32'd96;
end
262172:begin
	ram_in<=32'd96;
end
262173:begin
	ram_in<=32'd224;
end
262174:begin
	ram_in<=32'd96;
end
262175:begin
	ram_in<=32'd96;
end
262400:begin
	ram_in<=32'd76;
end
262401:begin
	ram_in<=32'd76;
end
262402:begin
	ram_in<=32'd236;
end
262403:begin
	ram_in<=32'd508;
end
262404:begin
	ram_in<=32'd476;
end
262405:begin
	ram_in<=32'd988;
end
262406:begin
	ram_in<=32'd984;
end
262407:begin
	ram_in<=32'd920;
end
262408:begin
	ram_in<=32'd1816;
end
262409:begin
	ram_in<=32'd3640;
end
262410:begin
	ram_in<=32'd3640;
end
262411:begin
	ram_in<=32'd3640;
end
262412:begin
	ram_in<=32'd3640;
end
262413:begin
	ram_in<=32'd7224;
end
262414:begin
	ram_in<=32'd7544;
end
262415:begin
	ram_in<=32'd8184;
end
262416:begin
	ram_in<=32'd8188;
end
262417:begin
	ram_in<=32'd8188;
end
262418:begin
	ram_in<=32'd8188;
end
262419:begin
	ram_in<=32'd8184;
end
262420:begin
	ram_in<=32'd4080;
end
262421:begin
	ram_in<=32'd96;
end
262422:begin
	ram_in<=32'd96;
end
262423:begin
	ram_in<=32'd96;
end
262424:begin
	ram_in<=32'd96;
end
262425:begin
	ram_in<=32'd192;
end
262426:begin
	ram_in<=32'd192;
end
262427:begin
	ram_in<=32'd192;
end
262428:begin
	ram_in<=32'd192;
end
262429:begin
	ram_in<=32'd192;
end
262430:begin
	ram_in<=32'd192;
end
262431:begin
	ram_in<=32'd192;
end
262656:begin
	ram_in<=32'd96;
end
262657:begin
	ram_in<=32'd112;
end
262658:begin
	ram_in<=32'd248;
end
262659:begin
	ram_in<=32'd248;
end
262660:begin
	ram_in<=32'd492;
end
262661:begin
	ram_in<=32'd508;
end
262662:begin
	ram_in<=32'd1944;
end
262663:begin
	ram_in<=32'd3992;
end
262664:begin
	ram_in<=32'd3864;
end
262665:begin
	ram_in<=32'd3608;
end
262666:begin
	ram_in<=32'd7704;
end
262667:begin
	ram_in<=32'd8184;
end
262668:begin
	ram_in<=32'd8184;
end
262669:begin
	ram_in<=32'd8184;
end
262670:begin
	ram_in<=32'd8188;
end
262671:begin
	ram_in<=32'd4092;
end
262672:begin
	ram_in<=32'd4092;
end
262673:begin
	ram_in<=32'd56;
end
262674:begin
	ram_in<=32'd48;
end
262675:begin
	ram_in<=32'd48;
end
262676:begin
	ram_in<=32'd96;
end
262677:begin
	ram_in<=32'd96;
end
262678:begin
	ram_in<=32'd96;
end
262679:begin
	ram_in<=32'd96;
end
262680:begin
	ram_in<=32'd96;
end
262681:begin
	ram_in<=32'd96;
end
262682:begin
	ram_in<=32'd96;
end
262683:begin
	ram_in<=32'd224;
end
262684:begin
	ram_in<=32'd224;
end
262685:begin
	ram_in<=32'd224;
end
262686:begin
	ram_in<=32'd224;
end
262687:begin
	ram_in<=32'd96;
end
262912:begin
	ram_in<=32'd96;
end
262913:begin
	ram_in<=32'd192;
end
262914:begin
	ram_in<=32'd192;
end
262915:begin
	ram_in<=32'd224;
end
262916:begin
	ram_in<=32'd192;
end
262917:begin
	ram_in<=32'd384;
end
262918:begin
	ram_in<=32'd896;
end
262919:begin
	ram_in<=32'd896;
end
262920:begin
	ram_in<=32'd896;
end
262921:begin
	ram_in<=32'd896;
end
262922:begin
	ram_in<=32'd1792;
end
262923:begin
	ram_in<=32'd1808;
end
262924:begin
	ram_in<=32'd1560;
end
262925:begin
	ram_in<=32'd1560;
end
262926:begin
	ram_in<=32'd3632;
end
262927:begin
	ram_in<=32'd3640;
end
262928:begin
	ram_in<=32'd3120;
end
262929:begin
	ram_in<=32'd3120;
end
262930:begin
	ram_in<=32'd3184;
end
262931:begin
	ram_in<=32'd7416;
end
262932:begin
	ram_in<=32'd8184;
end
262933:begin
	ram_in<=32'd8184;
end
262934:begin
	ram_in<=32'd8184;
end
262935:begin
	ram_in<=32'd8176;
end
262936:begin
	ram_in<=32'd4064;
end
262937:begin
	ram_in<=32'd224;
end
262938:begin
	ram_in<=32'd224;
end
262939:begin
	ram_in<=32'd224;
end
262940:begin
	ram_in<=32'd224;
end
262941:begin
	ram_in<=32'd224;
end
262942:begin
	ram_in<=32'd224;
end
262943:begin
	ram_in<=32'd96;
end
263168:begin
	ram_in<=32'd64;
end
263169:begin
	ram_in<=32'd224;
end
263170:begin
	ram_in<=32'd224;
end
263171:begin
	ram_in<=32'd192;
end
263172:begin
	ram_in<=32'd448;
end
263173:begin
	ram_in<=32'd448;
end
263174:begin
	ram_in<=32'd448;
end
263175:begin
	ram_in<=32'd448;
end
263176:begin
	ram_in<=32'd896;
end
263177:begin
	ram_in<=32'd904;
end
263178:begin
	ram_in<=32'd920;
end
263179:begin
	ram_in<=32'd924;
end
263180:begin
	ram_in<=32'd924;
end
263181:begin
	ram_in<=32'd1820;
end
263182:begin
	ram_in<=32'd3896;
end
263183:begin
	ram_in<=32'd3640;
end
263184:begin
	ram_in<=32'd3640;
end
263185:begin
	ram_in<=32'd3644;
end
263186:begin
	ram_in<=32'd8188;
end
263187:begin
	ram_in<=32'd8184;
end
263188:begin
	ram_in<=32'd16376;
end
263189:begin
	ram_in<=32'd16376;
end
263190:begin
	ram_in<=32'd16376;
end
263191:begin
	ram_in<=32'd8176;
end
263192:begin
	ram_in<=32'd8176;
end
263193:begin
	ram_in<=32'd224;
end
263194:begin
	ram_in<=32'd224;
end
263195:begin
	ram_in<=32'd224;
end
263196:begin
	ram_in<=32'd224;
end
263197:begin
	ram_in<=32'd240;
end
263198:begin
	ram_in<=32'd224;
end
263199:begin
	ram_in<=32'd224;
end
263424:begin
	ram_in<=32'd64;
end
263425:begin
	ram_in<=32'd192;
end
263426:begin
	ram_in<=32'd448;
end
263427:begin
	ram_in<=32'd448;
end
263428:begin
	ram_in<=32'd448;
end
263429:begin
	ram_in<=32'd448;
end
263430:begin
	ram_in<=32'd384;
end
263431:begin
	ram_in<=32'd896;
end
263432:begin
	ram_in<=32'd896;
end
263433:begin
	ram_in<=32'd896;
end
263434:begin
	ram_in<=32'd1800;
end
263435:begin
	ram_in<=32'd1800;
end
263436:begin
	ram_in<=32'd1560;
end
263437:begin
	ram_in<=32'd3612;
end
263438:begin
	ram_in<=32'd3612;
end
263439:begin
	ram_in<=32'd3096;
end
263440:begin
	ram_in<=32'd7224;
end
263441:begin
	ram_in<=32'd7224;
end
263442:begin
	ram_in<=32'd8176;
end
263443:begin
	ram_in<=32'd8176;
end
263444:begin
	ram_in<=32'd8176;
end
263445:begin
	ram_in<=32'd4080;
end
263446:begin
	ram_in<=32'd4080;
end
263447:begin
	ram_in<=32'd224;
end
263448:begin
	ram_in<=32'd224;
end
263449:begin
	ram_in<=32'd224;
end
263450:begin
	ram_in<=32'd224;
end
263451:begin
	ram_in<=32'd224;
end
263452:begin
	ram_in<=32'd224;
end
263453:begin
	ram_in<=32'd448;
end
263454:begin
	ram_in<=32'd224;
end
263455:begin
	ram_in<=32'd192;
end
263680:begin
	ram_in<=32'd96;
end
263681:begin
	ram_in<=32'd224;
end
263682:begin
	ram_in<=32'd480;
end
263683:begin
	ram_in<=32'd480;
end
263684:begin
	ram_in<=32'd480;
end
263685:begin
	ram_in<=32'd960;
end
263686:begin
	ram_in<=32'd896;
end
263687:begin
	ram_in<=32'd896;
end
263688:begin
	ram_in<=32'd1920;
end
263689:begin
	ram_in<=32'd1792;
end
263690:begin
	ram_in<=32'd1804;
end
263691:begin
	ram_in<=32'd3612;
end
263692:begin
	ram_in<=32'd3612;
end
263693:begin
	ram_in<=32'd3612;
end
263694:begin
	ram_in<=32'd3612;
end
263695:begin
	ram_in<=32'd7228;
end
263696:begin
	ram_in<=32'd7228;
end
263697:begin
	ram_in<=32'd7224;
end
263698:begin
	ram_in<=32'd15480;
end
263699:begin
	ram_in<=32'd7280;
end
263700:begin
	ram_in<=32'd8176;
end
263701:begin
	ram_in<=32'd8176;
end
263702:begin
	ram_in<=32'd16368;
end
263703:begin
	ram_in<=32'd8184;
end
263704:begin
	ram_in<=32'd4080;
end
263705:begin
	ram_in<=32'd4064;
end
263706:begin
	ram_in<=32'd480;
end
263707:begin
	ram_in<=32'd224;
end
263708:begin
	ram_in<=32'd480;
end
263709:begin
	ram_in<=32'd480;
end
263710:begin
	ram_in<=32'd480;
end
263711:begin
	ram_in<=32'd192;
end
263936:begin
	ram_in<=32'd128;
end
263937:begin
	ram_in<=32'd192;
end
263938:begin
	ram_in<=32'd192;
end
263939:begin
	ram_in<=32'd448;
end
263940:begin
	ram_in<=32'd448;
end
263941:begin
	ram_in<=32'd384;
end
263942:begin
	ram_in<=32'd896;
end
263943:begin
	ram_in<=32'd768;
end
263944:begin
	ram_in<=32'd768;
end
263945:begin
	ram_in<=32'd1792;
end
263946:begin
	ram_in<=32'd1792;
end
263947:begin
	ram_in<=32'd1808;
end
263948:begin
	ram_in<=32'd3632;
end
263949:begin
	ram_in<=32'd3632;
end
263950:begin
	ram_in<=32'd3632;
end
263951:begin
	ram_in<=32'd3184;
end
263952:begin
	ram_in<=32'd3184;
end
263953:begin
	ram_in<=32'd7216;
end
263954:begin
	ram_in<=32'd7264;
end
263955:begin
	ram_in<=32'd7264;
end
263956:begin
	ram_in<=32'd7280;
end
263957:begin
	ram_in<=32'd8176;
end
263958:begin
	ram_in<=32'd8176;
end
263959:begin
	ram_in<=32'd8176;
end
263960:begin
	ram_in<=32'd8160;
end
263961:begin
	ram_in<=32'd4032;
end
263962:begin
	ram_in<=32'd448;
end
263963:begin
	ram_in<=32'd448;
end
263964:begin
	ram_in<=32'd192;
end
263965:begin
	ram_in<=32'd192;
end
263966:begin
	ram_in<=32'd448;
end
263967:begin
	ram_in<=32'd128;
end
264192:begin
	ram_in<=32'd96;
end
264193:begin
	ram_in<=32'd96;
end
264194:begin
	ram_in<=32'd96;
end
264195:begin
	ram_in<=32'd192;
end
264196:begin
	ram_in<=32'd192;
end
264197:begin
	ram_in<=32'd192;
end
264198:begin
	ram_in<=32'd192;
end
264199:begin
	ram_in<=32'd448;
end
264200:begin
	ram_in<=32'd448;
end
264201:begin
	ram_in<=32'd448;
end
264202:begin
	ram_in<=32'd384;
end
264203:begin
	ram_in<=32'd384;
end
264204:begin
	ram_in<=32'd776;
end
264205:begin
	ram_in<=32'd780;
end
264206:begin
	ram_in<=32'd780;
end
264207:begin
	ram_in<=32'd1816;
end
264208:begin
	ram_in<=32'd1560;
end
264209:begin
	ram_in<=32'd1560;
end
264210:begin
	ram_in<=32'd3128;
end
264211:begin
	ram_in<=32'd3128;
end
264212:begin
	ram_in<=32'd7608;
end
264213:begin
	ram_in<=32'd8176;
end
264214:begin
	ram_in<=32'd8176;
end
264215:begin
	ram_in<=32'd8176;
end
264216:begin
	ram_in<=32'd8176;
end
264217:begin
	ram_in<=32'd8176;
end
264218:begin
	ram_in<=32'd6240;
end
264219:begin
	ram_in<=32'd96;
end
264220:begin
	ram_in<=32'd96;
end
264221:begin
	ram_in<=32'd96;
end
264222:begin
	ram_in<=32'd192;
end
264223:begin
	ram_in<=32'd64;
end
264448:begin
	ram_in<=32'd192;
end
264449:begin
	ram_in<=32'd448;
end
264450:begin
	ram_in<=32'd448;
end
264451:begin
	ram_in<=32'd448;
end
264452:begin
	ram_in<=32'd448;
end
264453:begin
	ram_in<=32'd960;
end
264454:begin
	ram_in<=32'd448;
end
264455:begin
	ram_in<=32'd896;
end
264456:begin
	ram_in<=32'd896;
end
264457:begin
	ram_in<=32'd896;
end
264458:begin
	ram_in<=32'd904;
end
264459:begin
	ram_in<=32'd1816;
end
264460:begin
	ram_in<=32'd1820;
end
264461:begin
	ram_in<=32'd3640;
end
264462:begin
	ram_in<=32'd3640;
end
264463:begin
	ram_in<=32'd3640;
end
264464:begin
	ram_in<=32'd3640;
end
264465:begin
	ram_in<=32'd7224;
end
264466:begin
	ram_in<=32'd7664;
end
264467:begin
	ram_in<=32'd16376;
end
264468:begin
	ram_in<=32'd16368;
end
264469:begin
	ram_in<=32'd16376;
end
264470:begin
	ram_in<=32'd16368;
end
264471:begin
	ram_in<=32'd16368;
end
264472:begin
	ram_in<=32'd16352;
end
264473:begin
	ram_in<=32'd6624;
end
264474:begin
	ram_in<=32'd448;
end
264475:begin
	ram_in<=32'd448;
end
264476:begin
	ram_in<=32'd448;
end
264477:begin
	ram_in<=32'd448;
end
264478:begin
	ram_in<=32'd448;
end
264479:begin
	ram_in<=32'd384;
end
327680:begin
	ram_in<=32'd352;
end
327681:begin
	ram_in<=32'd1016;
end
327682:begin
	ram_in<=32'd2044;
end
327683:begin
	ram_in<=32'd2044;
end
327684:begin
	ram_in<=32'd1924;
end
327685:begin
	ram_in<=32'd1792;
end
327686:begin
	ram_in<=32'd3072;
end
327687:begin
	ram_in<=32'd3072;
end
327688:begin
	ram_in<=32'd3264;
end
327689:begin
	ram_in<=32'd3264;
end
327690:begin
	ram_in<=32'd4080;
end
327691:begin
	ram_in<=32'd4080;
end
327692:begin
	ram_in<=32'd4088;
end
327693:begin
	ram_in<=32'd4080;
end
327694:begin
	ram_in<=32'd3960;
end
327695:begin
	ram_in<=32'd3640;
end
327696:begin
	ram_in<=32'd3128;
end
327697:begin
	ram_in<=32'd3128;
end
327698:begin
	ram_in<=32'd24;
end
327699:begin
	ram_in<=32'd24;
end
327700:begin
	ram_in<=32'd24;
end
327701:begin
	ram_in<=32'd24;
end
327702:begin
	ram_in<=32'd56;
end
327703:begin
	ram_in<=32'd48;
end
327704:begin
	ram_in<=32'd1584;
end
327705:begin
	ram_in<=32'd1648;
end
327706:begin
	ram_in<=32'd2032;
end
327707:begin
	ram_in<=32'd2016;
end
327708:begin
	ram_in<=32'd1984;
end
327709:begin
	ram_in<=32'd1984;
end
327710:begin
	ram_in<=32'd1920;
end
327711:begin
	ram_in<=32'd512;
end
327936:begin
	ram_in<=32'd32;
end
327937:begin
	ram_in<=32'd248;
end
327938:begin
	ram_in<=32'd504;
end
327939:begin
	ram_in<=32'd1016;
end
327940:begin
	ram_in<=32'd1984;
end
327941:begin
	ram_in<=32'd3968;
end
327942:begin
	ram_in<=32'd3840;
end
327943:begin
	ram_in<=32'd3584;
end
327944:begin
	ram_in<=32'd3584;
end
327945:begin
	ram_in<=32'd3584;
end
327946:begin
	ram_in<=32'd3072;
end
327947:begin
	ram_in<=32'd3072;
end
327948:begin
	ram_in<=32'd3168;
end
327949:begin
	ram_in<=32'd3312;
end
327950:begin
	ram_in<=32'd4080;
end
327951:begin
	ram_in<=32'd8184;
end
327952:begin
	ram_in<=32'd8088;
end
327953:begin
	ram_in<=32'd7960;
end
327954:begin
	ram_in<=32'd7704;
end
327955:begin
	ram_in<=32'd3096;
end
327956:begin
	ram_in<=32'd24;
end
327957:begin
	ram_in<=32'd24;
end
327958:begin
	ram_in<=32'd24;
end
327959:begin
	ram_in<=32'd56;
end
327960:begin
	ram_in<=32'd48;
end
327961:begin
	ram_in<=32'd48;
end
327962:begin
	ram_in<=32'd368;
end
327963:begin
	ram_in<=32'd480;
end
327964:begin
	ram_in<=32'd480;
end
327965:begin
	ram_in<=32'd480;
end
327966:begin
	ram_in<=32'd192;
end
327967:begin
	ram_in<=32'd128;
end
328192:begin
	ram_in<=32'd824;
end
328193:begin
	ram_in<=32'd1020;
end
328194:begin
	ram_in<=32'd1020;
end
328195:begin
	ram_in<=32'd2044;
end
328196:begin
	ram_in<=32'd2040;
end
328197:begin
	ram_in<=32'd1920;
end
328198:begin
	ram_in<=32'd1536;
end
328199:begin
	ram_in<=32'd1536;
end
328200:begin
	ram_in<=32'd3072;
end
328201:begin
	ram_in<=32'd3072;
end
328202:begin
	ram_in<=32'd3312;
end
328203:begin
	ram_in<=32'd3320;
end
328204:begin
	ram_in<=32'd8184;
end
328205:begin
	ram_in<=32'd8184;
end
328206:begin
	ram_in<=32'd8088;
end
328207:begin
	ram_in<=32'd7704;
end
328208:begin
	ram_in<=32'd3096;
end
328209:begin
	ram_in<=32'd24;
end
328210:begin
	ram_in<=32'd24;
end
328211:begin
	ram_in<=32'd24;
end
328212:begin
	ram_in<=32'd24;
end
328213:begin
	ram_in<=32'd48;
end
328214:begin
	ram_in<=32'd112;
end
328215:begin
	ram_in<=32'd96;
end
328216:begin
	ram_in<=32'd96;
end
328217:begin
	ram_in<=32'd96;
end
328218:begin
	ram_in<=32'd736;
end
328219:begin
	ram_in<=32'd960;
end
328220:begin
	ram_in<=32'd1984;
end
328221:begin
	ram_in<=32'd896;
end
328222:begin
	ram_in<=32'd1792;
end
328223:begin
	ram_in<=32'd768;
end
328448:begin
	ram_in<=32'd960;
end
328449:begin
	ram_in<=32'd1008;
end
328450:begin
	ram_in<=32'd2044;
end
328451:begin
	ram_in<=32'd2040;
end
328452:begin
	ram_in<=32'd2044;
end
328453:begin
	ram_in<=32'd4088;
end
328454:begin
	ram_in<=32'd3584;
end
328455:begin
	ram_in<=32'd1536;
end
328456:begin
	ram_in<=32'd3584;
end
328457:begin
	ram_in<=32'd3072;
end
328458:begin
	ram_in<=32'd3168;
end
328459:begin
	ram_in<=32'd3312;
end
328460:begin
	ram_in<=32'd7664;
end
328461:begin
	ram_in<=32'd8184;
end
328462:begin
	ram_in<=32'd8184;
end
328463:begin
	ram_in<=32'd8184;
end
328464:begin
	ram_in<=32'd7960;
end
328465:begin
	ram_in<=32'd7704;
end
328466:begin
	ram_in<=32'd7192;
end
328467:begin
	ram_in<=32'd7192;
end
328468:begin
	ram_in<=32'd24;
end
328469:begin
	ram_in<=32'd48;
end
328470:begin
	ram_in<=32'd48;
end
328471:begin
	ram_in<=32'd48;
end
328472:begin
	ram_in<=32'd112;
end
328473:begin
	ram_in<=32'd1632;
end
328474:begin
	ram_in<=32'd1760;
end
328475:begin
	ram_in<=32'd2016;
end
328476:begin
	ram_in<=32'd1984;
end
328477:begin
	ram_in<=32'd1984;
end
328478:begin
	ram_in<=32'd1920;
end
328479:begin
	ram_in<=32'd768;
end
328704:begin
	ram_in<=32'd16;
end
328705:begin
	ram_in<=32'd120;
end
328706:begin
	ram_in<=32'd2552;
end
328707:begin
	ram_in<=32'd4088;
end
328708:begin
	ram_in<=32'd4088;
end
328709:begin
	ram_in<=32'd4088;
end
328710:begin
	ram_in<=32'd4080;
end
328711:begin
	ram_in<=32'd3584;
end
328712:begin
	ram_in<=32'd3584;
end
328713:begin
	ram_in<=32'd3072;
end
328714:begin
	ram_in<=32'd3072;
end
328715:begin
	ram_in<=32'd3072;
end
328716:begin
	ram_in<=32'd4032;
end
328717:begin
	ram_in<=32'd4032;
end
328718:begin
	ram_in<=32'd8160;
end
328719:begin
	ram_in<=32'd8160;
end
328720:begin
	ram_in<=32'd8160;
end
328721:begin
	ram_in<=32'd3168;
end
328722:begin
	ram_in<=32'd96;
end
328723:begin
	ram_in<=32'd112;
end
328724:begin
	ram_in<=32'd112;
end
328725:begin
	ram_in<=32'd112;
end
328726:begin
	ram_in<=32'd112;
end
328727:begin
	ram_in<=32'd96;
end
328728:begin
	ram_in<=32'd224;
end
328729:begin
	ram_in<=32'd224;
end
328730:begin
	ram_in<=32'd960;
end
328731:begin
	ram_in<=32'd960;
end
328732:begin
	ram_in<=32'd3968;
end
328733:begin
	ram_in<=32'd3840;
end
328734:begin
	ram_in<=32'd3840;
end
328735:begin
	ram_in<=32'd3584;
end
328960:begin
	ram_in<=32'd0;
end
328961:begin
	ram_in<=32'd248;
end
328962:begin
	ram_in<=32'd2044;
end
328963:begin
	ram_in<=32'd4092;
end
328964:begin
	ram_in<=32'd4092;
end
328965:begin
	ram_in<=32'd4092;
end
328966:begin
	ram_in<=32'd3584;
end
328967:begin
	ram_in<=32'd3584;
end
328968:begin
	ram_in<=32'd3584;
end
328969:begin
	ram_in<=32'd3584;
end
328970:begin
	ram_in<=32'd1536;
end
328971:begin
	ram_in<=32'd4032;
end
328972:begin
	ram_in<=32'd4064;
end
328973:begin
	ram_in<=32'd2032;
end
328974:begin
	ram_in<=32'd2032;
end
328975:begin
	ram_in<=32'd4088;
end
328976:begin
	ram_in<=32'd2040;
end
328977:begin
	ram_in<=32'd1848;
end
328978:begin
	ram_in<=32'd1080;
end
328979:begin
	ram_in<=32'd56;
end
328980:begin
	ram_in<=32'd56;
end
328981:begin
	ram_in<=32'd56;
end
328982:begin
	ram_in<=32'd56;
end
328983:begin
	ram_in<=32'd112;
end
328984:begin
	ram_in<=32'd112;
end
328985:begin
	ram_in<=32'd240;
end
328986:begin
	ram_in<=32'd224;
end
328987:begin
	ram_in<=32'd992;
end
328988:begin
	ram_in<=32'd1984;
end
328989:begin
	ram_in<=32'd4032;
end
328990:begin
	ram_in<=32'd3968;
end
328991:begin
	ram_in<=32'd3840;
end
329216:begin
	ram_in<=32'd16;
end
329217:begin
	ram_in<=32'd368;
end
329218:begin
	ram_in<=32'd2040;
end
329219:begin
	ram_in<=32'd2040;
end
329220:begin
	ram_in<=32'd2040;
end
329221:begin
	ram_in<=32'd2040;
end
329222:begin
	ram_in<=32'd2032;
end
329223:begin
	ram_in<=32'd1792;
end
329224:begin
	ram_in<=32'd1536;
end
329225:begin
	ram_in<=32'd1536;
end
329226:begin
	ram_in<=32'd3584;
end
329227:begin
	ram_in<=32'd3584;
end
329228:begin
	ram_in<=32'd3072;
end
329229:begin
	ram_in<=32'd3072;
end
329230:begin
	ram_in<=32'd8176;
end
329231:begin
	ram_in<=32'd4080;
end
329232:begin
	ram_in<=32'd4088;
end
329233:begin
	ram_in<=32'd4088;
end
329234:begin
	ram_in<=32'd4088;
end
329235:begin
	ram_in<=32'd56;
end
329236:begin
	ram_in<=32'd24;
end
329237:begin
	ram_in<=32'd24;
end
329238:begin
	ram_in<=32'd24;
end
329239:begin
	ram_in<=32'd56;
end
329240:begin
	ram_in<=32'd48;
end
329241:begin
	ram_in<=32'd240;
end
329242:begin
	ram_in<=32'd496;
end
329243:begin
	ram_in<=32'd992;
end
329244:begin
	ram_in<=32'd2016;
end
329245:begin
	ram_in<=32'd1984;
end
329246:begin
	ram_in<=32'd1920;
end
329247:begin
	ram_in<=32'd1024;
end
329472:begin
	ram_in<=32'd24;
end
329473:begin
	ram_in<=32'd1016;
end
329474:begin
	ram_in<=32'd4088;
end
329475:begin
	ram_in<=32'd4088;
end
329476:begin
	ram_in<=32'd4088;
end
329477:begin
	ram_in<=32'd4064;
end
329478:begin
	ram_in<=32'd3840;
end
329479:begin
	ram_in<=32'd3584;
end
329480:begin
	ram_in<=32'd3072;
end
329481:begin
	ram_in<=32'd3072;
end
329482:begin
	ram_in<=32'd3072;
end
329483:begin
	ram_in<=32'd3072;
end
329484:begin
	ram_in<=32'd7168;
end
329485:begin
	ram_in<=32'd7680;
end
329486:begin
	ram_in<=32'd3968;
end
329487:begin
	ram_in<=32'd8128;
end
329488:begin
	ram_in<=32'd4032;
end
329489:begin
	ram_in<=32'd2016;
end
329490:begin
	ram_in<=32'd992;
end
329491:begin
	ram_in<=32'd112;
end
329492:begin
	ram_in<=32'd112;
end
329493:begin
	ram_in<=32'd112;
end
329494:begin
	ram_in<=32'd112;
end
329495:begin
	ram_in<=32'd112;
end
329496:begin
	ram_in<=32'd224;
end
329497:begin
	ram_in<=32'd2528;
end
329498:begin
	ram_in<=32'd3552;
end
329499:begin
	ram_in<=32'd4032;
end
329500:begin
	ram_in<=32'd4032;
end
329501:begin
	ram_in<=32'd3968;
end
329502:begin
	ram_in<=32'd3968;
end
329503:begin
	ram_in<=32'd1536;
end
329728:begin
	ram_in<=32'd128;
end
329729:begin
	ram_in<=32'd992;
end
329730:begin
	ram_in<=32'd2032;
end
329731:begin
	ram_in<=32'd2032;
end
329732:begin
	ram_in<=32'd2032;
end
329733:begin
	ram_in<=32'd2032;
end
329734:begin
	ram_in<=32'd1792;
end
329735:begin
	ram_in<=32'd3584;
end
329736:begin
	ram_in<=32'd3584;
end
329737:begin
	ram_in<=32'd3072;
end
329738:begin
	ram_in<=32'd3072;
end
329739:begin
	ram_in<=32'd3072;
end
329740:begin
	ram_in<=32'd3072;
end
329741:begin
	ram_in<=32'd8160;
end
329742:begin
	ram_in<=32'd4080;
end
329743:begin
	ram_in<=32'd4080;
end
329744:begin
	ram_in<=32'd4080;
end
329745:begin
	ram_in<=32'd4080;
end
329746:begin
	ram_in<=32'd48;
end
329747:begin
	ram_in<=32'd24;
end
329748:begin
	ram_in<=32'd24;
end
329749:begin
	ram_in<=32'd24;
end
329750:begin
	ram_in<=32'd56;
end
329751:begin
	ram_in<=32'd24;
end
329752:begin
	ram_in<=32'd120;
end
329753:begin
	ram_in<=32'd112;
end
329754:begin
	ram_in<=32'd240;
end
329755:begin
	ram_in<=32'd4064;
end
329756:begin
	ram_in<=32'd2016;
end
329757:begin
	ram_in<=32'd2016;
end
329758:begin
	ram_in<=32'd1984;
end
329759:begin
	ram_in<=32'd512;
end
329984:begin
	ram_in<=32'd896;
end
329985:begin
	ram_in<=32'd2016;
end
329986:begin
	ram_in<=32'd4080;
end
329987:begin
	ram_in<=32'd4080;
end
329988:begin
	ram_in<=32'd4080;
end
329989:begin
	ram_in<=32'd4088;
end
329990:begin
	ram_in<=32'd4088;
end
329991:begin
	ram_in<=32'd3864;
end
329992:begin
	ram_in<=32'd3856;
end
329993:begin
	ram_in<=32'd3584;
end
329994:begin
	ram_in<=32'd3840;
end
329995:begin
	ram_in<=32'd3584;
end
329996:begin
	ram_in<=32'd3584;
end
329997:begin
	ram_in<=32'd7680;
end
329998:begin
	ram_in<=32'd3584;
end
329999:begin
	ram_in<=32'd3968;
end
330000:begin
	ram_in<=32'd4032;
end
330001:begin
	ram_in<=32'd4032;
end
330002:begin
	ram_in<=32'd4064;
end
330003:begin
	ram_in<=32'd2016;
end
330004:begin
	ram_in<=32'd2032;
end
330005:begin
	ram_in<=32'd240;
end
330006:begin
	ram_in<=32'd96;
end
330007:begin
	ram_in<=32'd112;
end
330008:begin
	ram_in<=32'd112;
end
330009:begin
	ram_in<=32'd240;
end
330010:begin
	ram_in<=32'd2032;
end
330011:begin
	ram_in<=32'd4064;
end
330012:begin
	ram_in<=32'd4064;
end
330013:begin
	ram_in<=32'd4064;
end
330014:begin
	ram_in<=32'd2016;
end
330015:begin
	ram_in<=32'd1984;
end
393216:begin
	ram_in<=32'd256;
end
393217:begin
	ram_in<=32'd384;
end
393218:begin
	ram_in<=32'd448;
end
393219:begin
	ram_in<=32'd960;
end
393220:begin
	ram_in<=32'd896;
end
393221:begin
	ram_in<=32'd960;
end
393222:begin
	ram_in<=32'd960;
end
393223:begin
	ram_in<=32'd1792;
end
393224:begin
	ram_in<=32'd1792;
end
393225:begin
	ram_in<=32'd1792;
end
393226:begin
	ram_in<=32'd3840;
end
393227:begin
	ram_in<=32'd3584;
end
393228:begin
	ram_in<=32'd3584;
end
393229:begin
	ram_in<=32'd3584;
end
393230:begin
	ram_in<=32'd3584;
end
393231:begin
	ram_in<=32'd3808;
end
393232:begin
	ram_in<=32'd4080;
end
393233:begin
	ram_in<=32'd4080;
end
393234:begin
	ram_in<=32'd4088;
end
393235:begin
	ram_in<=32'd4024;
end
393236:begin
	ram_in<=32'd3596;
end
393237:begin
	ram_in<=32'd3596;
end
393238:begin
	ram_in<=32'd3596;
end
393239:begin
	ram_in<=32'd1542;
end
393240:begin
	ram_in<=32'd1542;
end
393241:begin
	ram_in<=32'd1798;
end
393242:begin
	ram_in<=32'd1822;
end
393243:begin
	ram_in<=32'd1854;
end
393244:begin
	ram_in<=32'd1020;
end
393245:begin
	ram_in<=32'd508;
end
393246:begin
	ram_in<=32'd508;
end
393247:begin
	ram_in<=32'd240;
end
393472:begin
	ram_in<=32'd256;
end
393473:begin
	ram_in<=32'd256;
end
393474:begin
	ram_in<=32'd896;
end
393475:begin
	ram_in<=32'd960;
end
393476:begin
	ram_in<=32'd960;
end
393477:begin
	ram_in<=32'd1920;
end
393478:begin
	ram_in<=32'd960;
end
393479:begin
	ram_in<=32'd1920;
end
393480:begin
	ram_in<=32'd1792;
end
393481:begin
	ram_in<=32'd1792;
end
393482:begin
	ram_in<=32'd3840;
end
393483:begin
	ram_in<=32'd3584;
end
393484:begin
	ram_in<=32'd1536;
end
393485:begin
	ram_in<=32'd1536;
end
393486:begin
	ram_in<=32'd3584;
end
393487:begin
	ram_in<=32'd1536;
end
393488:begin
	ram_in<=32'd4032;
end
393489:begin
	ram_in<=32'd4064;
end
393490:begin
	ram_in<=32'd2032;
end
393491:begin
	ram_in<=32'd2040;
end
393492:begin
	ram_in<=32'd2040;
end
393493:begin
	ram_in<=32'd1820;
end
393494:begin
	ram_in<=32'd1564;
end
393495:begin
	ram_in<=32'd1548;
end
393496:begin
	ram_in<=32'd1806;
end
393497:begin
	ram_in<=32'd798;
end
393498:begin
	ram_in<=32'd828;
end
393499:begin
	ram_in<=32'd1022;
end
393500:begin
	ram_in<=32'd1020;
end
393501:begin
	ram_in<=32'd1020;
end
393502:begin
	ram_in<=32'd248;
end
393503:begin
	ram_in<=32'd224;
end
393728:begin
	ram_in<=32'd128;
end
393729:begin
	ram_in<=32'd448;
end
393730:begin
	ram_in<=32'd960;
end
393731:begin
	ram_in<=32'd992;
end
393732:begin
	ram_in<=32'd992;
end
393733:begin
	ram_in<=32'd1984;
end
393734:begin
	ram_in<=32'd1920;
end
393735:begin
	ram_in<=32'd1920;
end
393736:begin
	ram_in<=32'd1792;
end
393737:begin
	ram_in<=32'd1792;
end
393738:begin
	ram_in<=32'd1792;
end
393739:begin
	ram_in<=32'd1792;
end
393740:begin
	ram_in<=32'd1536;
end
393741:begin
	ram_in<=32'd1536;
end
393742:begin
	ram_in<=32'd3584;
end
393743:begin
	ram_in<=32'd2016;
end
393744:begin
	ram_in<=32'd2016;
end
393745:begin
	ram_in<=32'd2032;
end
393746:begin
	ram_in<=32'd2040;
end
393747:begin
	ram_in<=32'd4088;
end
393748:begin
	ram_in<=32'd4092;
end
393749:begin
	ram_in<=32'd3964;
end
393750:begin
	ram_in<=32'd3854;
end
393751:begin
	ram_in<=32'd3854;
end
393752:begin
	ram_in<=32'd3870;
end
393753:begin
	ram_in<=32'd3868;
end
393754:begin
	ram_in<=32'd2044;
end
393755:begin
	ram_in<=32'd2044;
end
393756:begin
	ram_in<=32'd1016;
end
393757:begin
	ram_in<=32'd1016;
end
393758:begin
	ram_in<=32'd496;
end
393759:begin
	ram_in<=32'd480;
end
393984:begin
	ram_in<=32'd192;
end
393985:begin
	ram_in<=32'd224;
end
393986:begin
	ram_in<=32'd1008;
end
393987:begin
	ram_in<=32'd1008;
end
393988:begin
	ram_in<=32'd1008;
end
393989:begin
	ram_in<=32'd1008;
end
393990:begin
	ram_in<=32'd1920;
end
393991:begin
	ram_in<=32'd1792;
end
393992:begin
	ram_in<=32'd1536;
end
393993:begin
	ram_in<=32'd3584;
end
393994:begin
	ram_in<=32'd1536;
end
393995:begin
	ram_in<=32'd3584;
end
393996:begin
	ram_in<=32'd3584;
end
393997:begin
	ram_in<=32'd3168;
end
393998:begin
	ram_in<=32'd3824;
end
393999:begin
	ram_in<=32'd4080;
end
394000:begin
	ram_in<=32'd4088;
end
394001:begin
	ram_in<=32'd4088;
end
394002:begin
	ram_in<=32'd4024;
end
394003:begin
	ram_in<=32'd3996;
end
394004:begin
	ram_in<=32'd3868;
end
394005:begin
	ram_in<=32'd3596;
end
394006:begin
	ram_in<=32'd3596;
end
394007:begin
	ram_in<=32'd1548;
end
394008:begin
	ram_in<=32'd1804;
end
394009:begin
	ram_in<=32'd1820;
end
394010:begin
	ram_in<=32'd1980;
end
394011:begin
	ram_in<=32'd2044;
end
394012:begin
	ram_in<=32'd1020;
end
394013:begin
	ram_in<=32'd1020;
end
394014:begin
	ram_in<=32'd504;
end
394015:begin
	ram_in<=32'd96;
end
394240:begin
	ram_in<=32'd256;
end
394241:begin
	ram_in<=32'd896;
end
394242:begin
	ram_in<=32'd896;
end
394243:begin
	ram_in<=32'd896;
end
394244:begin
	ram_in<=32'd1920;
end
394245:begin
	ram_in<=32'd1920;
end
394246:begin
	ram_in<=32'd1792;
end
394247:begin
	ram_in<=32'd1792;
end
394248:begin
	ram_in<=32'd1536;
end
394249:begin
	ram_in<=32'd1536;
end
394250:begin
	ram_in<=32'd1536;
end
394251:begin
	ram_in<=32'd1536;
end
394252:begin
	ram_in<=32'd3584;
end
394253:begin
	ram_in<=32'd3072;
end
394254:begin
	ram_in<=32'd3584;
end
394255:begin
	ram_in<=32'd3584;
end
394256:begin
	ram_in<=32'd4064;
end
394257:begin
	ram_in<=32'd4080;
end
394258:begin
	ram_in<=32'd4088;
end
394259:begin
	ram_in<=32'd4092;
end
394260:begin
	ram_in<=32'd4092;
end
394261:begin
	ram_in<=32'd3596;
end
394262:begin
	ram_in<=32'd3084;
end
394263:begin
	ram_in<=32'd3596;
end
394264:begin
	ram_in<=32'd1548;
end
394265:begin
	ram_in<=32'd1548;
end
394266:begin
	ram_in<=32'd1548;
end
394267:begin
	ram_in<=32'd1820;
end
394268:begin
	ram_in<=32'd956;
end
394269:begin
	ram_in<=32'd1016;
end
394270:begin
	ram_in<=32'd504;
end
394271:begin
	ram_in<=32'd240;
end
394496:begin
	ram_in<=32'd192;
end
394497:begin
	ram_in<=32'd448;
end
394498:begin
	ram_in<=32'd992;
end
394499:begin
	ram_in<=32'd960;
end
394500:begin
	ram_in<=32'd1984;
end
394501:begin
	ram_in<=32'd1920;
end
394502:begin
	ram_in<=32'd1920;
end
394503:begin
	ram_in<=32'd1792;
end
394504:begin
	ram_in<=32'd3840;
end
394505:begin
	ram_in<=32'd3584;
end
394506:begin
	ram_in<=32'd3584;
end
394507:begin
	ram_in<=32'd3072;
end
394508:begin
	ram_in<=32'd6144;
end
394509:begin
	ram_in<=32'd2048;
end
394510:begin
	ram_in<=32'd2112;
end
394511:begin
	ram_in<=32'd6256;
end
394512:begin
	ram_in<=32'd6256;
end
394513:begin
	ram_in<=32'd6256;
end
394514:begin
	ram_in<=32'd6264;
end
394515:begin
	ram_in<=32'd8184;
end
394516:begin
	ram_in<=32'd3608;
end
394517:begin
	ram_in<=32'd3612;
end
394518:begin
	ram_in<=32'd3612;
end
394519:begin
	ram_in<=32'd3608;
end
394520:begin
	ram_in<=32'd3608;
end
394521:begin
	ram_in<=32'd3608;
end
394522:begin
	ram_in<=32'd1976;
end
394523:begin
	ram_in<=32'd2044;
end
394524:begin
	ram_in<=32'd1016;
end
394525:begin
	ram_in<=32'd1016;
end
394526:begin
	ram_in<=32'd504;
end
394527:begin
	ram_in<=32'd32;
end
394752:begin
	ram_in<=32'd128;
end
394753:begin
	ram_in<=32'd192;
end
394754:begin
	ram_in<=32'd448;
end
394755:begin
	ram_in<=32'd448;
end
394756:begin
	ram_in<=32'd960;
end
394757:begin
	ram_in<=32'd960;
end
394758:begin
	ram_in<=32'd896;
end
394759:begin
	ram_in<=32'd1920;
end
394760:begin
	ram_in<=32'd896;
end
394761:begin
	ram_in<=32'd768;
end
394762:begin
	ram_in<=32'd1792;
end
394763:begin
	ram_in<=32'd1792;
end
394764:begin
	ram_in<=32'd1536;
end
394765:begin
	ram_in<=32'd1792;
end
394766:begin
	ram_in<=32'd1792;
end
394767:begin
	ram_in<=32'd1536;
end
394768:begin
	ram_in<=32'd1536;
end
394769:begin
	ram_in<=32'd3584;
end
394770:begin
	ram_in<=32'd1792;
end
394771:begin
	ram_in<=32'd3968;
end
394772:begin
	ram_in<=32'd4088;
end
394773:begin
	ram_in<=32'd4088;
end
394774:begin
	ram_in<=32'd4092;
end
394775:begin
	ram_in<=32'd1918;
end
394776:begin
	ram_in<=32'd1566;
end
394777:begin
	ram_in<=32'd1806;
end
394778:begin
	ram_in<=32'd1934;
end
394779:begin
	ram_in<=32'd958;
end
394780:begin
	ram_in<=32'd510;
end
394781:begin
	ram_in<=32'd510;
end
394782:begin
	ram_in<=32'd508;
end
394783:begin
	ram_in<=32'd112;
end
395008:begin
	ram_in<=32'd128;
end
395009:begin
	ram_in<=32'd960;
end
395010:begin
	ram_in<=32'd960;
end
395011:begin
	ram_in<=32'd960;
end
395012:begin
	ram_in<=32'd896;
end
395013:begin
	ram_in<=32'd1792;
end
395014:begin
	ram_in<=32'd1792;
end
395015:begin
	ram_in<=32'd1792;
end
395016:begin
	ram_in<=32'd1536;
end
395017:begin
	ram_in<=32'd1536;
end
395018:begin
	ram_in<=32'd1536;
end
395019:begin
	ram_in<=32'd1536;
end
395020:begin
	ram_in<=32'd1536;
end
395021:begin
	ram_in<=32'd3584;
end
395022:begin
	ram_in<=32'd3584;
end
395023:begin
	ram_in<=32'd1536;
end
395024:begin
	ram_in<=32'd1536;
end
395025:begin
	ram_in<=32'd3584;
end
395026:begin
	ram_in<=32'd3824;
end
395027:begin
	ram_in<=32'd4088;
end
395028:begin
	ram_in<=32'd4088;
end
395029:begin
	ram_in<=32'd4092;
end
395030:begin
	ram_in<=32'd2044;
end
395031:begin
	ram_in<=32'd1804;
end
395032:begin
	ram_in<=32'd1548;
end
395033:begin
	ram_in<=32'd1548;
end
395034:begin
	ram_in<=32'd1804;
end
395035:begin
	ram_in<=32'd2044;
end
395036:begin
	ram_in<=32'd2044;
end
395037:begin
	ram_in<=32'd1016;
end
395038:begin
	ram_in<=32'd504;
end
395039:begin
	ram_in<=32'd64;
end
395264:begin
	ram_in<=32'd384;
end
395265:begin
	ram_in<=32'd448;
end
395266:begin
	ram_in<=32'd960;
end
395267:begin
	ram_in<=32'd896;
end
395268:begin
	ram_in<=32'd896;
end
395269:begin
	ram_in<=32'd1920;
end
395270:begin
	ram_in<=32'd896;
end
395271:begin
	ram_in<=32'd1792;
end
395272:begin
	ram_in<=32'd1792;
end
395273:begin
	ram_in<=32'd1792;
end
395274:begin
	ram_in<=32'd1792;
end
395275:begin
	ram_in<=32'd1536;
end
395276:begin
	ram_in<=32'd3584;
end
395277:begin
	ram_in<=32'd1792;
end
395278:begin
	ram_in<=32'd1792;
end
395279:begin
	ram_in<=32'd3584;
end
395280:begin
	ram_in<=32'd3584;
end
395281:begin
	ram_in<=32'd4080;
end
395282:begin
	ram_in<=32'd4088;
end
395283:begin
	ram_in<=32'd4088;
end
395284:begin
	ram_in<=32'd4092;
end
395285:begin
	ram_in<=32'd4092;
end
395286:begin
	ram_in<=32'd8188;
end
395287:begin
	ram_in<=32'd3596;
end
395288:begin
	ram_in<=32'd3852;
end
395289:begin
	ram_in<=32'd1804;
end
395290:begin
	ram_in<=32'd1820;
end
395291:begin
	ram_in<=32'd1022;
end
395292:begin
	ram_in<=32'd1020;
end
395293:begin
	ram_in<=32'd1020;
end
395294:begin
	ram_in<=32'd508;
end
395295:begin
	ram_in<=32'd248;
end
395520:begin
	ram_in<=32'd512;
end
395521:begin
	ram_in<=32'd768;
end
395522:begin
	ram_in<=32'd768;
end
395523:begin
	ram_in<=32'd768;
end
395524:begin
	ram_in<=32'd1792;
end
395525:begin
	ram_in<=32'd1792;
end
395526:begin
	ram_in<=32'd1536;
end
395527:begin
	ram_in<=32'd3584;
end
395528:begin
	ram_in<=32'd3584;
end
395529:begin
	ram_in<=32'd3072;
end
395530:begin
	ram_in<=32'd7168;
end
395531:begin
	ram_in<=32'd6144;
end
395532:begin
	ram_in<=32'd3072;
end
395533:begin
	ram_in<=32'd3072;
end
395534:begin
	ram_in<=32'd2048;
end
395535:begin
	ram_in<=32'd2048;
end
395536:begin
	ram_in<=32'd2048;
end
395537:begin
	ram_in<=32'd6256;
end
395538:begin
	ram_in<=32'd2296;
end
395539:begin
	ram_in<=32'd3576;
end
395540:begin
	ram_in<=32'd4088;
end
395541:begin
	ram_in<=32'd4092;
end
395542:begin
	ram_in<=32'd4092;
end
395543:begin
	ram_in<=32'd4060;
end
395544:begin
	ram_in<=32'd1820;
end
395545:begin
	ram_in<=32'd1852;
end
395546:begin
	ram_in<=32'd1912;
end
395547:begin
	ram_in<=32'd2032;
end
395548:begin
	ram_in<=32'd2032;
end
395549:begin
	ram_in<=32'd992;
end
395550:begin
	ram_in<=32'd992;
end
395551:begin
	ram_in<=32'd384;
end
458752:begin
	ram_in<=32'd63;
end
458753:begin
	ram_in<=32'd127;
end
458754:begin
	ram_in<=32'd1023;
end
458755:begin
	ram_in<=32'd2047;
end
458756:begin
	ram_in<=32'd2047;
end
458757:begin
	ram_in<=32'd2046;
end
458758:begin
	ram_in<=32'd1934;
end
458759:begin
	ram_in<=32'd1822;
end
458760:begin
	ram_in<=32'd28;
end
458761:begin
	ram_in<=32'd24;
end
458762:begin
	ram_in<=32'd56;
end
458763:begin
	ram_in<=32'd56;
end
458764:begin
	ram_in<=32'd48;
end
458765:begin
	ram_in<=32'd112;
end
458766:begin
	ram_in<=32'd1016;
end
458767:begin
	ram_in<=32'd2040;
end
458768:begin
	ram_in<=32'd2044;
end
458769:begin
	ram_in<=32'd2040;
end
458770:begin
	ram_in<=32'd4080;
end
458771:begin
	ram_in<=32'd2016;
end
458772:begin
	ram_in<=32'd224;
end
458773:begin
	ram_in<=32'd192;
end
458774:begin
	ram_in<=32'd448;
end
458775:begin
	ram_in<=32'd192;
end
458776:begin
	ram_in<=32'd448;
end
458777:begin
	ram_in<=32'd448;
end
458778:begin
	ram_in<=32'd448;
end
458779:begin
	ram_in<=32'd896;
end
458780:begin
	ram_in<=32'd896;
end
458781:begin
	ram_in<=32'd896;
end
458782:begin
	ram_in<=32'd896;
end
458783:begin
	ram_in<=32'd256;
end
459008:begin
	ram_in<=32'd48;
end
459009:begin
	ram_in<=32'd504;
end
459010:begin
	ram_in<=32'd1020;
end
459011:begin
	ram_in<=32'd2044;
end
459012:begin
	ram_in<=32'd2044;
end
459013:begin
	ram_in<=32'd2044;
end
459014:begin
	ram_in<=32'd1564;
end
459015:begin
	ram_in<=32'd1052;
end
459016:begin
	ram_in<=32'd28;
end
459017:begin
	ram_in<=32'd28;
end
459018:begin
	ram_in<=32'd24;
end
459019:begin
	ram_in<=32'd24;
end
459020:begin
	ram_in<=32'd24;
end
459021:begin
	ram_in<=32'd4088;
end
459022:begin
	ram_in<=32'd8184;
end
459023:begin
	ram_in<=32'd8184;
end
459024:begin
	ram_in<=32'd8184;
end
459025:begin
	ram_in<=32'd8176;
end
459026:begin
	ram_in<=32'd3936;
end
459027:begin
	ram_in<=32'd224;
end
459028:begin
	ram_in<=32'd224;
end
459029:begin
	ram_in<=32'd224;
end
459030:begin
	ram_in<=32'd224;
end
459031:begin
	ram_in<=32'd448;
end
459032:begin
	ram_in<=32'd448;
end
459033:begin
	ram_in<=32'd384;
end
459034:begin
	ram_in<=32'd384;
end
459035:begin
	ram_in<=32'd896;
end
459036:begin
	ram_in<=32'd896;
end
459037:begin
	ram_in<=32'd896;
end
459038:begin
	ram_in<=32'd768;
end
459039:begin
	ram_in<=32'd768;
end
459264:begin
	ram_in<=32'd248;
end
459265:begin
	ram_in<=32'd1020;
end
459266:begin
	ram_in<=32'd2044;
end
459267:begin
	ram_in<=32'd2044;
end
459268:begin
	ram_in<=32'd2046;
end
459269:begin
	ram_in<=32'd2046;
end
459270:begin
	ram_in<=32'd3868;
end
459271:begin
	ram_in<=32'd1052;
end
459272:begin
	ram_in<=32'd28;
end
459273:begin
	ram_in<=32'd56;
end
459274:begin
	ram_in<=32'd632;
end
459275:begin
	ram_in<=32'd1020;
end
459276:begin
	ram_in<=32'd2044;
end
459277:begin
	ram_in<=32'd2044;
end
459278:begin
	ram_in<=32'd2044;
end
459279:begin
	ram_in<=32'd4088;
end
459280:begin
	ram_in<=32'd2016;
end
459281:begin
	ram_in<=32'd224;
end
459282:begin
	ram_in<=32'd448;
end
459283:begin
	ram_in<=32'd448;
end
459284:begin
	ram_in<=32'd448;
end
459285:begin
	ram_in<=32'd448;
end
459286:begin
	ram_in<=32'd448;
end
459287:begin
	ram_in<=32'd448;
end
459288:begin
	ram_in<=32'd896;
end
459289:begin
	ram_in<=32'd896;
end
459290:begin
	ram_in<=32'd896;
end
459291:begin
	ram_in<=32'd1920;
end
459292:begin
	ram_in<=32'd1920;
end
459293:begin
	ram_in<=32'd1920;
end
459294:begin
	ram_in<=32'd1792;
end
459295:begin
	ram_in<=32'd1792;
end
459520:begin
	ram_in<=32'd240;
end
459521:begin
	ram_in<=32'd504;
end
459522:begin
	ram_in<=32'd1016;
end
459523:begin
	ram_in<=32'd2040;
end
459524:begin
	ram_in<=32'd2044;
end
459525:begin
	ram_in<=32'd1564;
end
459526:begin
	ram_in<=32'd3096;
end
459527:begin
	ram_in<=32'd24;
end
459528:begin
	ram_in<=32'd24;
end
459529:begin
	ram_in<=32'd24;
end
459530:begin
	ram_in<=32'd56;
end
459531:begin
	ram_in<=32'd56;
end
459532:begin
	ram_in<=32'd56;
end
459533:begin
	ram_in<=32'd3824;
end
459534:begin
	ram_in<=32'd8184;
end
459535:begin
	ram_in<=32'd8184;
end
459536:begin
	ram_in<=32'd8176;
end
459537:begin
	ram_in<=32'd3808;
end
459538:begin
	ram_in<=32'd224;
end
459539:begin
	ram_in<=32'd224;
end
459540:begin
	ram_in<=32'd192;
end
459541:begin
	ram_in<=32'd192;
end
459542:begin
	ram_in<=32'd384;
end
459543:begin
	ram_in<=32'd384;
end
459544:begin
	ram_in<=32'd384;
end
459545:begin
	ram_in<=32'd384;
end
459546:begin
	ram_in<=32'd384;
end
459547:begin
	ram_in<=32'd768;
end
459548:begin
	ram_in<=32'd768;
end
459549:begin
	ram_in<=32'd768;
end
459550:begin
	ram_in<=32'd896;
end
459551:begin
	ram_in<=32'd768;
end
459776:begin
	ram_in<=32'd120;
end
459777:begin
	ram_in<=32'd2040;
end
459778:begin
	ram_in<=32'd2044;
end
459779:begin
	ram_in<=32'd4088;
end
459780:begin
	ram_in<=32'd4092;
end
459781:begin
	ram_in<=32'd4092;
end
459782:begin
	ram_in<=32'd1948;
end
459783:begin
	ram_in<=32'd1048;
end
459784:begin
	ram_in<=32'd56;
end
459785:begin
	ram_in<=32'd56;
end
459786:begin
	ram_in<=32'd48;
end
459787:begin
	ram_in<=32'd48;
end
459788:begin
	ram_in<=32'd112;
end
459789:begin
	ram_in<=32'd1144;
end
459790:begin
	ram_in<=32'd4088;
end
459791:begin
	ram_in<=32'd4092;
end
459792:begin
	ram_in<=32'd4092;
end
459793:begin
	ram_in<=32'd4092;
end
459794:begin
	ram_in<=32'd4092;
end
459795:begin
	ram_in<=32'd4088;
end
459796:begin
	ram_in<=32'd2008;
end
459797:begin
	ram_in<=32'd400;
end
459798:begin
	ram_in<=32'd384;
end
459799:begin
	ram_in<=32'd896;
end
459800:begin
	ram_in<=32'd896;
end
459801:begin
	ram_in<=32'd768;
end
459802:begin
	ram_in<=32'd1792;
end
459803:begin
	ram_in<=32'd1792;
end
459804:begin
	ram_in<=32'd1792;
end
459805:begin
	ram_in<=32'd1792;
end
459806:begin
	ram_in<=32'd1536;
end
459807:begin
	ram_in<=32'd1536;
end
460032:begin
	ram_in<=32'd960;
end
460033:begin
	ram_in<=32'd2016;
end
460034:begin
	ram_in<=32'd4080;
end
460035:begin
	ram_in<=32'd4080;
end
460036:begin
	ram_in<=32'd4088;
end
460037:begin
	ram_in<=32'd1080;
end
460038:begin
	ram_in<=32'd56;
end
460039:begin
	ram_in<=32'd24;
end
460040:begin
	ram_in<=32'd56;
end
460041:begin
	ram_in<=32'd56;
end
460042:begin
	ram_in<=32'd48;
end
460043:begin
	ram_in<=32'd112;
end
460044:begin
	ram_in<=32'd112;
end
460045:begin
	ram_in<=32'd96;
end
460046:begin
	ram_in<=32'd96;
end
460047:begin
	ram_in<=32'd3296;
end
460048:begin
	ram_in<=32'd4088;
end
460049:begin
	ram_in<=32'd4088;
end
460050:begin
	ram_in<=32'd4088;
end
460051:begin
	ram_in<=32'd4088;
end
460052:begin
	ram_in<=32'd960;
end
460053:begin
	ram_in<=32'd384;
end
460054:begin
	ram_in<=32'd384;
end
460055:begin
	ram_in<=32'd768;
end
460056:begin
	ram_in<=32'd768;
end
460057:begin
	ram_in<=32'd1792;
end
460058:begin
	ram_in<=32'd1792;
end
460059:begin
	ram_in<=32'd1792;
end
460060:begin
	ram_in<=32'd1536;
end
460061:begin
	ram_in<=32'd3584;
end
460062:begin
	ram_in<=32'd1536;
end
460063:begin
	ram_in<=32'd1536;
end
460288:begin
	ram_in<=32'd28;
end
460289:begin
	ram_in<=32'd510;
end
460290:begin
	ram_in<=32'd1022;
end
460291:begin
	ram_in<=32'd2046;
end
460292:begin
	ram_in<=32'd4094;
end
460293:begin
	ram_in<=32'd4094;
end
460294:begin
	ram_in<=32'd2046;
end
460295:begin
	ram_in<=32'd3598;
end
460296:begin
	ram_in<=32'd1038;
end
460297:begin
	ram_in<=32'd30;
end
460298:begin
	ram_in<=32'd28;
end
460299:begin
	ram_in<=32'd28;
end
460300:begin
	ram_in<=32'd28;
end
460301:begin
	ram_in<=32'd280;
end
460302:begin
	ram_in<=32'd504;
end
460303:begin
	ram_in<=32'd1016;
end
460304:begin
	ram_in<=32'd1016;
end
460305:begin
	ram_in<=32'd1016;
end
460306:begin
	ram_in<=32'd2032;
end
460307:begin
	ram_in<=32'd1008;
end
460308:begin
	ram_in<=32'd1008;
end
460309:begin
	ram_in<=32'd224;
end
460310:begin
	ram_in<=32'd192;
end
460311:begin
	ram_in<=32'd448;
end
460312:begin
	ram_in<=32'd448;
end
460313:begin
	ram_in<=32'd448;
end
460314:begin
	ram_in<=32'd960;
end
460315:begin
	ram_in<=32'd960;
end
460316:begin
	ram_in<=32'd896;
end
460317:begin
	ram_in<=32'd896;
end
460318:begin
	ram_in<=32'd896;
end
460319:begin
	ram_in<=32'd768;
end
460544:begin
	ram_in<=32'd992;
end
460545:begin
	ram_in<=32'd1008;
end
460546:begin
	ram_in<=32'd2032;
end
460547:begin
	ram_in<=32'd4080;
end
460548:begin
	ram_in<=32'd4080;
end
460549:begin
	ram_in<=32'd4088;
end
460550:begin
	ram_in<=32'd1912;
end
460551:begin
	ram_in<=32'd1080;
end
460552:begin
	ram_in<=32'd56;
end
460553:begin
	ram_in<=32'd56;
end
460554:begin
	ram_in<=32'd56;
end
460555:begin
	ram_in<=32'd112;
end
460556:begin
	ram_in<=32'd112;
end
460557:begin
	ram_in<=32'd112;
end
460558:begin
	ram_in<=32'd112;
end
460559:begin
	ram_in<=32'd112;
end
460560:begin
	ram_in<=32'd1008;
end
460561:begin
	ram_in<=32'd2032;
end
460562:begin
	ram_in<=32'd4088;
end
460563:begin
	ram_in<=32'd4088;
end
460564:begin
	ram_in<=32'd4088;
end
460565:begin
	ram_in<=32'd4088;
end
460566:begin
	ram_in<=32'd4080;
end
460567:begin
	ram_in<=32'd960;
end
460568:begin
	ram_in<=32'd960;
end
460569:begin
	ram_in<=32'd896;
end
460570:begin
	ram_in<=32'd896;
end
460571:begin
	ram_in<=32'd1920;
end
460572:begin
	ram_in<=32'd1792;
end
460573:begin
	ram_in<=32'd1792;
end
460574:begin
	ram_in<=32'd1792;
end
460575:begin
	ram_in<=32'd1536;
end
460800:begin
	ram_in<=32'd504;
end
460801:begin
	ram_in<=32'd1016;
end
460802:begin
	ram_in<=32'd2040;
end
460803:begin
	ram_in<=32'd2044;
end
460804:begin
	ram_in<=32'd4092;
end
460805:begin
	ram_in<=32'd4092;
end
460806:begin
	ram_in<=32'd3644;
end
460807:begin
	ram_in<=32'd3612;
end
460808:begin
	ram_in<=32'd1052;
end
460809:begin
	ram_in<=32'd28;
end
460810:begin
	ram_in<=32'd60;
end
460811:begin
	ram_in<=32'd56;
end
460812:begin
	ram_in<=32'd56;
end
460813:begin
	ram_in<=32'd56;
end
460814:begin
	ram_in<=32'd1016;
end
460815:begin
	ram_in<=32'd2040;
end
460816:begin
	ram_in<=32'd4092;
end
460817:begin
	ram_in<=32'd4092;
end
460818:begin
	ram_in<=32'd4092;
end
460819:begin
	ram_in<=32'd4088;
end
460820:begin
	ram_in<=32'd3808;
end
460821:begin
	ram_in<=32'd1248;
end
460822:begin
	ram_in<=32'd224;
end
460823:begin
	ram_in<=32'd448;
end
460824:begin
	ram_in<=32'd384;
end
460825:begin
	ram_in<=32'd896;
end
460826:begin
	ram_in<=32'd896;
end
460827:begin
	ram_in<=32'd896;
end
460828:begin
	ram_in<=32'd1792;
end
460829:begin
	ram_in<=32'd1792;
end
460830:begin
	ram_in<=32'd1792;
end
460831:begin
	ram_in<=32'd1536;
end
461056:begin
	ram_in<=32'd1008;
end
461057:begin
	ram_in<=32'd1016;
end
461058:begin
	ram_in<=32'd2040;
end
461059:begin
	ram_in<=32'd2040;
end
461060:begin
	ram_in<=32'd2040;
end
461061:begin
	ram_in<=32'd1660;
end
461062:begin
	ram_in<=32'd1084;
end
461063:begin
	ram_in<=32'd60;
end
461064:begin
	ram_in<=32'd60;
end
461065:begin
	ram_in<=32'd56;
end
461066:begin
	ram_in<=32'd56;
end
461067:begin
	ram_in<=32'd56;
end
461068:begin
	ram_in<=32'd112;
end
461069:begin
	ram_in<=32'd112;
end
461070:begin
	ram_in<=32'd112;
end
461071:begin
	ram_in<=32'd112;
end
461072:begin
	ram_in<=32'd112;
end
461073:begin
	ram_in<=32'd240;
end
461074:begin
	ram_in<=32'd4088;
end
461075:begin
	ram_in<=32'd4088;
end
461076:begin
	ram_in<=32'd4088;
end
461077:begin
	ram_in<=32'd8184;
end
461078:begin
	ram_in<=32'd4088;
end
461079:begin
	ram_in<=32'd4080;
end
461080:begin
	ram_in<=32'd3008;
end
461081:begin
	ram_in<=32'd896;
end
461082:begin
	ram_in<=32'd896;
end
461083:begin
	ram_in<=32'd896;
end
461084:begin
	ram_in<=32'd896;
end
461085:begin
	ram_in<=32'd1920;
end
461086:begin
	ram_in<=32'd1792;
end
461087:begin
	ram_in<=32'd1792;
end
524288:begin
	ram_in<=32'd0;
end
524289:begin
	ram_in<=32'd1984;
end
524290:begin
	ram_in<=32'd1984;
end
524291:begin
	ram_in<=32'd4064;
end
524292:begin
	ram_in<=32'd3696;
end
524293:begin
	ram_in<=32'd3632;
end
524294:begin
	ram_in<=32'd7216;
end
524295:begin
	ram_in<=32'd3120;
end
524296:begin
	ram_in<=32'd7216;
end
524297:begin
	ram_in<=32'd7280;
end
524298:begin
	ram_in<=32'd7408;
end
524299:begin
	ram_in<=32'd8160;
end
524300:begin
	ram_in<=32'd8160;
end
524301:begin
	ram_in<=32'd8128;
end
524302:begin
	ram_in<=32'd4032;
end
524303:begin
	ram_in<=32'd2016;
end
524304:begin
	ram_in<=32'd2016;
end
524305:begin
	ram_in<=32'd2016;
end
524306:begin
	ram_in<=32'd1936;
end
524307:begin
	ram_in<=32'd1808;
end
524308:begin
	ram_in<=32'd1552;
end
524309:begin
	ram_in<=32'd1560;
end
524310:begin
	ram_in<=32'd1544;
end
524311:begin
	ram_in<=32'd1560;
end
524312:begin
	ram_in<=32'd1560;
end
524313:begin
	ram_in<=32'd1560;
end
524314:begin
	ram_in<=32'd1560;
end
524315:begin
	ram_in<=32'd2040;
end
524316:begin
	ram_in<=32'd2032;
end
524317:begin
	ram_in<=32'd2032;
end
524318:begin
	ram_in<=32'd1008;
end
524319:begin
	ram_in<=32'd0;
end
524544:begin
	ram_in<=32'd448;
end
524545:begin
	ram_in<=32'd2016;
end
524546:begin
	ram_in<=32'd2032;
end
524547:begin
	ram_in<=32'd3888;
end
524548:begin
	ram_in<=32'd3120;
end
524549:begin
	ram_in<=32'd7224;
end
524550:begin
	ram_in<=32'd7224;
end
524551:begin
	ram_in<=32'd6256;
end
524552:begin
	ram_in<=32'd6640;
end
524553:begin
	ram_in<=32'd8160;
end
524554:begin
	ram_in<=32'd8160;
end
524555:begin
	ram_in<=32'd8064;
end
524556:begin
	ram_in<=32'd3968;
end
524557:begin
	ram_in<=32'd1984;
end
524558:begin
	ram_in<=32'd1984;
end
524559:begin
	ram_in<=32'd4064;
end
524560:begin
	ram_in<=32'd3936;
end
524561:begin
	ram_in<=32'd3696;
end
524562:begin
	ram_in<=32'd3120;
end
524563:begin
	ram_in<=32'd3088;
end
524564:begin
	ram_in<=32'd3096;
end
524565:begin
	ram_in<=32'd3096;
end
524566:begin
	ram_in<=32'd3100;
end
524567:begin
	ram_in<=32'd3084;
end
524568:begin
	ram_in<=32'd3096;
end
524569:begin
	ram_in<=32'd3096;
end
524570:begin
	ram_in<=32'd3128;
end
524571:begin
	ram_in<=32'd3696;
end
524572:begin
	ram_in<=32'd4080;
end
524573:begin
	ram_in<=32'd2016;
end
524574:begin
	ram_in<=32'd992;
end
524575:begin
	ram_in<=32'd896;
end
524800:begin
	ram_in<=32'd112;
end
524801:begin
	ram_in<=32'd240;
end
524802:begin
	ram_in<=32'd504;
end
524803:begin
	ram_in<=32'd1016;
end
524804:begin
	ram_in<=32'd2040;
end
524805:begin
	ram_in<=32'd2040;
end
524806:begin
	ram_in<=32'd7736;
end
524807:begin
	ram_in<=32'd7224;
end
524808:begin
	ram_in<=32'd7224;
end
524809:begin
	ram_in<=32'd7224;
end
524810:begin
	ram_in<=32'd3640;
end
524811:begin
	ram_in<=32'd3952;
end
524812:begin
	ram_in<=32'd2032;
end
524813:begin
	ram_in<=32'd2016;
end
524814:begin
	ram_in<=32'd2016;
end
524815:begin
	ram_in<=32'd992;
end
524816:begin
	ram_in<=32'd1008;
end
524817:begin
	ram_in<=32'd1008;
end
524818:begin
	ram_in<=32'd1008;
end
524819:begin
	ram_in<=32'd880;
end
524820:begin
	ram_in<=32'd1848;
end
524821:begin
	ram_in<=32'd1848;
end
524822:begin
	ram_in<=32'd1592;
end
524823:begin
	ram_in<=32'd792;
end
524824:begin
	ram_in<=32'd1816;
end
524825:begin
	ram_in<=32'd1848;
end
524826:begin
	ram_in<=32'd824;
end
524827:begin
	ram_in<=32'd1008;
end
524828:begin
	ram_in<=32'd1008;
end
524829:begin
	ram_in<=32'd480;
end
524830:begin
	ram_in<=32'd480;
end
524831:begin
	ram_in<=32'd128;
end
525056:begin
	ram_in<=32'd256;
end
525057:begin
	ram_in<=32'd992;
end
525058:begin
	ram_in<=32'd992;
end
525059:begin
	ram_in<=32'd2040;
end
525060:begin
	ram_in<=32'd2040;
end
525061:begin
	ram_in<=32'd1848;
end
525062:begin
	ram_in<=32'd3640;
end
525063:begin
	ram_in<=32'd7224;
end
525064:begin
	ram_in<=32'd7224;
end
525065:begin
	ram_in<=32'd7280;
end
525066:begin
	ram_in<=32'd6256;
end
525067:begin
	ram_in<=32'd6256;
end
525068:begin
	ram_in<=32'd7792;
end
525069:begin
	ram_in<=32'd3808;
end
525070:begin
	ram_in<=32'd4064;
end
525071:begin
	ram_in<=32'd4032;
end
525072:begin
	ram_in<=32'd1984;
end
525073:begin
	ram_in<=32'd960;
end
525074:begin
	ram_in<=32'd992;
end
525075:begin
	ram_in<=32'd992;
end
525076:begin
	ram_in<=32'd880;
end
525077:begin
	ram_in<=32'd824;
end
525078:begin
	ram_in<=32'd824;
end
525079:begin
	ram_in<=32'd1848;
end
525080:begin
	ram_in<=32'd1592;
end
525081:begin
	ram_in<=32'd1592;
end
525082:begin
	ram_in<=32'd1656;
end
525083:begin
	ram_in<=32'd1784;
end
525084:begin
	ram_in<=32'd2032;
end
525085:begin
	ram_in<=32'd992;
end
525086:begin
	ram_in<=32'd992;
end
525087:begin
	ram_in<=32'd480;
end
525312:begin
	ram_in<=32'd96;
end
525313:begin
	ram_in<=32'd496;
end
525314:begin
	ram_in<=32'd496;
end
525315:begin
	ram_in<=32'd1016;
end
525316:begin
	ram_in<=32'd2040;
end
525317:begin
	ram_in<=32'd1976;
end
525318:begin
	ram_in<=32'd1848;
end
525319:begin
	ram_in<=32'd1592;
end
525320:begin
	ram_in<=32'd7216;
end
525321:begin
	ram_in<=32'd7280;
end
525322:begin
	ram_in<=32'd7280;
end
525323:begin
	ram_in<=32'd7792;
end
525324:begin
	ram_in<=32'd8032;
end
525325:begin
	ram_in<=32'd4064;
end
525326:begin
	ram_in<=32'd4032;
end
525327:begin
	ram_in<=32'd1984;
end
525328:begin
	ram_in<=32'd960;
end
525329:begin
	ram_in<=32'd448;
end
525330:begin
	ram_in<=32'd480;
end
525331:begin
	ram_in<=32'd480;
end
525332:begin
	ram_in<=32'd496;
end
525333:begin
	ram_in<=32'd368;
end
525334:begin
	ram_in<=32'd368;
end
525335:begin
	ram_in<=32'd312;
end
525336:begin
	ram_in<=32'd312;
end
525337:begin
	ram_in<=32'd312;
end
525338:begin
	ram_in<=32'd368;
end
525339:begin
	ram_in<=32'd496;
end
525340:begin
	ram_in<=32'd496;
end
525341:begin
	ram_in<=32'd480;
end
525342:begin
	ram_in<=32'd480;
end
525343:begin
	ram_in<=32'd192;
end
525568:begin
	ram_in<=32'd384;
end
525569:begin
	ram_in<=32'd992;
end
525570:begin
	ram_in<=32'd2032;
end
525571:begin
	ram_in<=32'd2032;
end
525572:begin
	ram_in<=32'd2032;
end
525573:begin
	ram_in<=32'd2032;
end
525574:begin
	ram_in<=32'd3640;
end
525575:begin
	ram_in<=32'd7736;
end
525576:begin
	ram_in<=32'd7224;
end
525577:begin
	ram_in<=32'd7224;
end
525578:begin
	ram_in<=32'd7224;
end
525579:begin
	ram_in<=32'd3640;
end
525580:begin
	ram_in<=32'd3696;
end
525581:begin
	ram_in<=32'd4080;
end
525582:begin
	ram_in<=32'd4080;
end
525583:begin
	ram_in<=32'd2016;
end
525584:begin
	ram_in<=32'd992;
end
525585:begin
	ram_in<=32'd480;
end
525586:begin
	ram_in<=32'd992;
end
525587:begin
	ram_in<=32'd1008;
end
525588:begin
	ram_in<=32'd1008;
end
525589:begin
	ram_in<=32'd1904;
end
525590:begin
	ram_in<=32'd1840;
end
525591:begin
	ram_in<=32'd1848;
end
525592:begin
	ram_in<=32'd1560;
end
525593:begin
	ram_in<=32'd1560;
end
525594:begin
	ram_in<=32'd1592;
end
525595:begin
	ram_in<=32'd1912;
end
525596:begin
	ram_in<=32'd2040;
end
525597:begin
	ram_in<=32'd2032;
end
525598:begin
	ram_in<=32'd1008;
end
525599:begin
	ram_in<=32'd960;
end
525824:begin
	ram_in<=32'd256;
end
525825:begin
	ram_in<=32'd896;
end
525826:begin
	ram_in<=32'd896;
end
525827:begin
	ram_in<=32'd1984;
end
525828:begin
	ram_in<=32'd1984;
end
525829:begin
	ram_in<=32'd1984;
end
525830:begin
	ram_in<=32'd1728;
end
525831:begin
	ram_in<=32'd3776;
end
525832:begin
	ram_in<=32'd3648;
end
525833:begin
	ram_in<=32'd3584;
end
525834:begin
	ram_in<=32'd1544;
end
525835:begin
	ram_in<=32'd1848;
end
525836:begin
	ram_in<=32'd1912;
end
525837:begin
	ram_in<=32'd2040;
end
525838:begin
	ram_in<=32'd2040;
end
525839:begin
	ram_in<=32'd2016;
end
525840:begin
	ram_in<=32'd1984;
end
525841:begin
	ram_in<=32'd1920;
end
525842:begin
	ram_in<=32'd4032;
end
525843:begin
	ram_in<=32'd4032;
end
525844:begin
	ram_in<=32'd8160;
end
525845:begin
	ram_in<=32'd7392;
end
525846:begin
	ram_in<=32'd7408;
end
525847:begin
	ram_in<=32'd3184;
end
525848:begin
	ram_in<=32'd3128;
end
525849:begin
	ram_in<=32'd3128;
end
525850:begin
	ram_in<=32'd3608;
end
525851:begin
	ram_in<=32'd1564;
end
525852:begin
	ram_in<=32'd2044;
end
525853:begin
	ram_in<=32'd1020;
end
525854:begin
	ram_in<=32'd504;
end
525855:begin
	ram_in<=32'd496;
end
526080:begin
	ram_in<=32'd384;
end
526081:begin
	ram_in<=32'd960;
end
526082:begin
	ram_in<=32'd2016;
end
526083:begin
	ram_in<=32'd4064;
end
526084:begin
	ram_in<=32'd4064;
end
526085:begin
	ram_in<=32'd3808;
end
526086:begin
	ram_in<=32'd3680;
end
526087:begin
	ram_in<=32'd3168;
end
526088:begin
	ram_in<=32'd3168;
end
526089:begin
	ram_in<=32'd3616;
end
526090:begin
	ram_in<=32'd3584;
end
526091:begin
	ram_in<=32'd3584;
end
526092:begin
	ram_in<=32'd1792;
end
526093:begin
	ram_in<=32'd1816;
end
526094:begin
	ram_in<=32'd1848;
end
526095:begin
	ram_in<=32'd1016;
end
526096:begin
	ram_in<=32'd1016;
end
526097:begin
	ram_in<=32'd1016;
end
526098:begin
	ram_in<=32'd1016;
end
526099:begin
	ram_in<=32'd2016;
end
526100:begin
	ram_in<=32'd2016;
end
526101:begin
	ram_in<=32'd4064;
end
526102:begin
	ram_in<=32'd4064;
end
526103:begin
	ram_in<=32'd7904;
end
526104:begin
	ram_in<=32'd7264;
end
526105:begin
	ram_in<=32'd7280;
end
526106:begin
	ram_in<=32'd7280;
end
526107:begin
	ram_in<=32'd3696;
end
526108:begin
	ram_in<=32'd4080;
end
526109:begin
	ram_in<=32'd2016;
end
526110:begin
	ram_in<=32'd1984;
end
526111:begin
	ram_in<=32'd896;
end
526336:begin
	ram_in<=32'd128;
end
526337:begin
	ram_in<=32'd992;
end
526338:begin
	ram_in<=32'd2016;
end
526339:begin
	ram_in<=32'd2032;
end
526340:begin
	ram_in<=32'd2032;
end
526341:begin
	ram_in<=32'd1648;
end
526342:begin
	ram_in<=32'd1648;
end
526343:begin
	ram_in<=32'd1648;
end
526344:begin
	ram_in<=32'd1648;
end
526345:begin
	ram_in<=32'd1120;
end
526346:begin
	ram_in<=32'd7264;
end
526347:begin
	ram_in<=32'd3680;
end
526348:begin
	ram_in<=32'd8160;
end
526349:begin
	ram_in<=32'd4032;
end
526350:begin
	ram_in<=32'd4032;
end
526351:begin
	ram_in<=32'd960;
end
526352:begin
	ram_in<=32'd480;
end
526353:begin
	ram_in<=32'd480;
end
526354:begin
	ram_in<=32'd504;
end
526355:begin
	ram_in<=32'd312;
end
526356:begin
	ram_in<=32'd824;
end
526357:begin
	ram_in<=32'd536;
end
526358:begin
	ram_in<=32'd780;
end
526359:begin
	ram_in<=32'd1548;
end
526360:begin
	ram_in<=32'd1548;
end
526361:begin
	ram_in<=32'd1548;
end
526362:begin
	ram_in<=32'd1564;
end
526363:begin
	ram_in<=32'd1660;
end
526364:begin
	ram_in<=32'd1656;
end
526365:begin
	ram_in<=32'd2032;
end
526366:begin
	ram_in<=32'd992;
end
526367:begin
	ram_in<=32'd992;
end
526592:begin
	ram_in<=32'd192;
end
526593:begin
	ram_in<=32'd1008;
end
526594:begin
	ram_in<=32'd2032;
end
526595:begin
	ram_in<=32'd2032;
end
526596:begin
	ram_in<=32'd2032;
end
526597:begin
	ram_in<=32'd1904;
end
526598:begin
	ram_in<=32'd1648;
end
526599:begin
	ram_in<=32'd3184;
end
526600:begin
	ram_in<=32'd3184;
end
526601:begin
	ram_in<=32'd3296;
end
526602:begin
	ram_in<=32'd7392;
end
526603:begin
	ram_in<=32'd8128;
end
526604:begin
	ram_in<=32'd8128;
end
526605:begin
	ram_in<=32'd3968;
end
526606:begin
	ram_in<=32'd3968;
end
526607:begin
	ram_in<=32'd1984;
end
526608:begin
	ram_in<=32'd2016;
end
526609:begin
	ram_in<=32'd2032;
end
526610:begin
	ram_in<=32'd2032;
end
526611:begin
	ram_in<=32'd1648;
end
526612:begin
	ram_in<=32'd1656;
end
526613:begin
	ram_in<=32'd1592;
end
526614:begin
	ram_in<=32'd1592;
end
526615:begin
	ram_in<=32'd1560;
end
526616:begin
	ram_in<=32'd1560;
end
526617:begin
	ram_in<=32'd1560;
end
526618:begin
	ram_in<=32'd1560;
end
526619:begin
	ram_in<=32'd1784;
end
526620:begin
	ram_in<=32'd2040;
end
526621:begin
	ram_in<=32'd2040;
end
526622:begin
	ram_in<=32'd2032;
end
526623:begin
	ram_in<=32'd480;
end
589824:begin
	ram_in<=32'd96;
end
589825:begin
	ram_in<=32'd112;
end
589826:begin
	ram_in<=32'd240;
end
589827:begin
	ram_in<=32'd504;
end
589828:begin
	ram_in<=32'd1016;
end
589829:begin
	ram_in<=32'd1022;
end
589830:begin
	ram_in<=32'd958;
end
589831:begin
	ram_in<=32'd1820;
end
589832:begin
	ram_in<=32'd1804;
end
589833:begin
	ram_in<=32'd1804;
end
589834:begin
	ram_in<=32'd3644;
end
589835:begin
	ram_in<=32'd3708;
end
589836:begin
	ram_in<=32'd3320;
end
589837:begin
	ram_in<=32'd4088;
end
589838:begin
	ram_in<=32'd4088;
end
589839:begin
	ram_in<=32'd4024;
end
589840:begin
	ram_in<=32'd3896;
end
589841:begin
	ram_in<=32'd3128;
end
589842:begin
	ram_in<=32'd48;
end
589843:begin
	ram_in<=32'd48;
end
589844:begin
	ram_in<=32'd48;
end
589845:begin
	ram_in<=32'd112;
end
589846:begin
	ram_in<=32'd112;
end
589847:begin
	ram_in<=32'd96;
end
589848:begin
	ram_in<=32'd96;
end
589849:begin
	ram_in<=32'd96;
end
589850:begin
	ram_in<=32'd224;
end
589851:begin
	ram_in<=32'd224;
end
589852:begin
	ram_in<=32'd224;
end
589853:begin
	ram_in<=32'd224;
end
589854:begin
	ram_in<=32'd192;
end
589855:begin
	ram_in<=32'd128;
end
590080:begin
	ram_in<=32'd32;
end
590081:begin
	ram_in<=32'd116;
end
590082:begin
	ram_in<=32'd246;
end
590083:begin
	ram_in<=32'd508;
end
590084:begin
	ram_in<=32'd508;
end
590085:begin
	ram_in<=32'd414;
end
590086:begin
	ram_in<=32'd798;
end
590087:begin
	ram_in<=32'd1596;
end
590088:begin
	ram_in<=32'd1596;
end
590089:begin
	ram_in<=32'd1052;
end
590090:begin
	ram_in<=32'd1052;
end
590091:begin
	ram_in<=32'd3096;
end
590092:begin
	ram_in<=32'd3096;
end
590093:begin
	ram_in<=32'd3128;
end
590094:begin
	ram_in<=32'd3184;
end
590095:begin
	ram_in<=32'd2544;
end
590096:begin
	ram_in<=32'd4016;
end
590097:begin
	ram_in<=32'd4016;
end
590098:begin
	ram_in<=32'd3872;
end
590099:begin
	ram_in<=32'd3104;
end
590100:begin
	ram_in<=32'd32;
end
590101:begin
	ram_in<=32'd96;
end
590102:begin
	ram_in<=32'd96;
end
590103:begin
	ram_in<=32'd96;
end
590104:begin
	ram_in<=32'd96;
end
590105:begin
	ram_in<=32'd224;
end
590106:begin
	ram_in<=32'd192;
end
590107:begin
	ram_in<=32'd192;
end
590108:begin
	ram_in<=32'd192;
end
590109:begin
	ram_in<=32'd224;
end
590110:begin
	ram_in<=32'd192;
end
590111:begin
	ram_in<=32'd64;
end
590336:begin
	ram_in<=32'd56;
end
590337:begin
	ram_in<=32'd60;
end
590338:begin
	ram_in<=32'd252;
end
590339:begin
	ram_in<=32'd252;
end
590340:begin
	ram_in<=32'd508;
end
590341:begin
	ram_in<=32'd460;
end
590342:begin
	ram_in<=32'd924;
end
590343:begin
	ram_in<=32'd782;
end
590344:begin
	ram_in<=32'd782;
end
590345:begin
	ram_in<=32'd1550;
end
590346:begin
	ram_in<=32'd1550;
end
590347:begin
	ram_in<=32'd3100;
end
590348:begin
	ram_in<=32'd3196;
end
590349:begin
	ram_in<=32'd3324;
end
590350:begin
	ram_in<=32'd4092;
end
590351:begin
	ram_in<=32'd4056;
end
590352:begin
	ram_in<=32'd3992;
end
590353:begin
	ram_in<=32'd3864;
end
590354:begin
	ram_in<=32'd3608;
end
590355:begin
	ram_in<=32'd24;
end
590356:begin
	ram_in<=32'd48;
end
590357:begin
	ram_in<=32'd48;
end
590358:begin
	ram_in<=32'd48;
end
590359:begin
	ram_in<=32'd48;
end
590360:begin
	ram_in<=32'd96;
end
590361:begin
	ram_in<=32'd96;
end
590362:begin
	ram_in<=32'd96;
end
590363:begin
	ram_in<=32'd96;
end
590364:begin
	ram_in<=32'd96;
end
590365:begin
	ram_in<=32'd192;
end
590366:begin
	ram_in<=32'd192;
end
590367:begin
	ram_in<=32'd128;
end
590592:begin
	ram_in<=32'd32;
end
590593:begin
	ram_in<=32'd240;
end
590594:begin
	ram_in<=32'd504;
end
590595:begin
	ram_in<=32'd1008;
end
590596:begin
	ram_in<=32'd2040;
end
590597:begin
	ram_in<=32'd3896;
end
590598:begin
	ram_in<=32'd3608;
end
590599:begin
	ram_in<=32'd3096;
end
590600:begin
	ram_in<=32'd3096;
end
590601:begin
	ram_in<=32'd3096;
end
590602:begin
	ram_in<=32'd6168;
end
590603:begin
	ram_in<=32'd6200;
end
590604:begin
	ram_in<=32'd6200;
end
590605:begin
	ram_in<=32'd7288;
end
590606:begin
	ram_in<=32'd7416;
end
590607:begin
	ram_in<=32'd4088;
end
590608:begin
	ram_in<=32'd4088;
end
590609:begin
	ram_in<=32'd4088;
end
590610:begin
	ram_in<=32'd1968;
end
590611:begin
	ram_in<=32'd48;
end
590612:begin
	ram_in<=32'd112;
end
590613:begin
	ram_in<=32'd112;
end
590614:begin
	ram_in<=32'd96;
end
590615:begin
	ram_in<=32'd96;
end
590616:begin
	ram_in<=32'd224;
end
590617:begin
	ram_in<=32'd192;
end
590618:begin
	ram_in<=32'd192;
end
590619:begin
	ram_in<=32'd448;
end
590620:begin
	ram_in<=32'd448;
end
590621:begin
	ram_in<=32'd384;
end
590622:begin
	ram_in<=32'd896;
end
590623:begin
	ram_in<=32'd384;
end
590848:begin
	ram_in<=32'd504;
end
590849:begin
	ram_in<=32'd1016;
end
590850:begin
	ram_in<=32'd1020;
end
590851:begin
	ram_in<=32'd1020;
end
590852:begin
	ram_in<=32'd2044;
end
590853:begin
	ram_in<=32'd1932;
end
590854:begin
	ram_in<=32'd3612;
end
590855:begin
	ram_in<=32'd3612;
end
590856:begin
	ram_in<=32'd3100;
end
590857:begin
	ram_in<=32'd3100;
end
590858:begin
	ram_in<=32'd3132;
end
590859:begin
	ram_in<=32'd3192;
end
590860:begin
	ram_in<=32'd3192;
end
590861:begin
	ram_in<=32'd7664;
end
590862:begin
	ram_in<=32'd7664;
end
590863:begin
	ram_in<=32'd4080;
end
590864:begin
	ram_in<=32'd4080;
end
590865:begin
	ram_in<=32'd4080;
end
590866:begin
	ram_in<=32'd2032;
end
590867:begin
	ram_in<=32'd1888;
end
590868:begin
	ram_in<=32'd192;
end
590869:begin
	ram_in<=32'd192;
end
590870:begin
	ram_in<=32'd192;
end
590871:begin
	ram_in<=32'd448;
end
590872:begin
	ram_in<=32'd448;
end
590873:begin
	ram_in<=32'd448;
end
590874:begin
	ram_in<=32'd960;
end
590875:begin
	ram_in<=32'd896;
end
590876:begin
	ram_in<=32'd896;
end
590877:begin
	ram_in<=32'd896;
end
590878:begin
	ram_in<=32'd896;
end
590879:begin
	ram_in<=32'd768;
end
591104:begin
	ram_in<=32'd224;
end
591105:begin
	ram_in<=32'd240;
end
591106:begin
	ram_in<=32'd1016;
end
591107:begin
	ram_in<=32'd1008;
end
591108:begin
	ram_in<=32'd2040;
end
591109:begin
	ram_in<=32'd1848;
end
591110:begin
	ram_in<=32'd3612;
end
591111:begin
	ram_in<=32'd3100;
end
591112:begin
	ram_in<=32'd3100;
end
591113:begin
	ram_in<=32'd3100;
end
591114:begin
	ram_in<=32'd3100;
end
591115:begin
	ram_in<=32'd3132;
end
591116:begin
	ram_in<=32'd3320;
end
591117:begin
	ram_in<=32'd4088;
end
591118:begin
	ram_in<=32'd4088;
end
591119:begin
	ram_in<=32'd2032;
end
591120:begin
	ram_in<=32'd2032;
end
591121:begin
	ram_in<=32'd944;
end
591122:begin
	ram_in<=32'd112;
end
591123:begin
	ram_in<=32'd96;
end
591124:begin
	ram_in<=32'd96;
end
591125:begin
	ram_in<=32'd192;
end
591126:begin
	ram_in<=32'd192;
end
591127:begin
	ram_in<=32'd448;
end
591128:begin
	ram_in<=32'd448;
end
591129:begin
	ram_in<=32'd384;
end
591130:begin
	ram_in<=32'd384;
end
591131:begin
	ram_in<=32'd896;
end
591132:begin
	ram_in<=32'd896;
end
591133:begin
	ram_in<=32'd896;
end
591134:begin
	ram_in<=32'd768;
end
591135:begin
	ram_in<=32'd768;
end
591360:begin
	ram_in<=32'd448;
end
591361:begin
	ram_in<=32'd1008;
end
591362:begin
	ram_in<=32'd1008;
end
591363:begin
	ram_in<=32'd2040;
end
591364:begin
	ram_in<=32'd2040;
end
591365:begin
	ram_in<=32'd3900;
end
591366:begin
	ram_in<=32'd3612;
end
591367:begin
	ram_in<=32'd3612;
end
591368:begin
	ram_in<=32'd3612;
end
591369:begin
	ram_in<=32'd3100;
end
591370:begin
	ram_in<=32'd3128;
end
591371:begin
	ram_in<=32'd3832;
end
591372:begin
	ram_in<=32'd4088;
end
591373:begin
	ram_in<=32'd4088;
end
591374:begin
	ram_in<=32'd2040;
end
591375:begin
	ram_in<=32'd2040;
end
591376:begin
	ram_in<=32'd56;
end
591377:begin
	ram_in<=32'd48;
end
591378:begin
	ram_in<=32'd112;
end
591379:begin
	ram_in<=32'd112;
end
591380:begin
	ram_in<=32'd112;
end
591381:begin
	ram_in<=32'd112;
end
591382:begin
	ram_in<=32'd224;
end
591383:begin
	ram_in<=32'd224;
end
591384:begin
	ram_in<=32'd448;
end
591385:begin
	ram_in<=32'd448;
end
591386:begin
	ram_in<=32'd960;
end
591387:begin
	ram_in<=32'd960;
end
591388:begin
	ram_in<=32'd1984;
end
591389:begin
	ram_in<=32'd896;
end
591390:begin
	ram_in<=32'd896;
end
591391:begin
	ram_in<=32'd896;
end
591616:begin
	ram_in<=32'd128;
end
591617:begin
	ram_in<=32'd448;
end
591618:begin
	ram_in<=32'd960;
end
591619:begin
	ram_in<=32'd1984;
end
591620:begin
	ram_in<=32'd4032;
end
591621:begin
	ram_in<=32'd4080;
end
591622:begin
	ram_in<=32'd3696;
end
591623:begin
	ram_in<=32'd3184;
end
591624:begin
	ram_in<=32'd3184;
end
591625:begin
	ram_in<=32'd6256;
end
591626:begin
	ram_in<=32'd6384;
end
591627:begin
	ram_in<=32'd8176;
end
591628:begin
	ram_in<=32'd4080;
end
591629:begin
	ram_in<=32'd4080;
end
591630:begin
	ram_in<=32'd4080;
end
591631:begin
	ram_in<=32'd560;
end
591632:begin
	ram_in<=32'd48;
end
591633:begin
	ram_in<=32'd16;
end
591634:begin
	ram_in<=32'd24;
end
591635:begin
	ram_in<=32'd24;
end
591636:begin
	ram_in<=32'd24;
end
591637:begin
	ram_in<=32'd24;
end
591638:begin
	ram_in<=32'd8;
end
591639:begin
	ram_in<=32'd8;
end
591640:begin
	ram_in<=32'd8;
end
591641:begin
	ram_in<=32'd8;
end
591642:begin
	ram_in<=32'd1560;
end
591643:begin
	ram_in<=32'd1560;
end
591644:begin
	ram_in<=32'd2040;
end
591645:begin
	ram_in<=32'd1016;
end
591646:begin
	ram_in<=32'd2032;
end
591647:begin
	ram_in<=32'd448;
end
591872:begin
	ram_in<=32'd480;
end
591873:begin
	ram_in<=32'd992;
end
591874:begin
	ram_in<=32'd992;
end
591875:begin
	ram_in<=32'd2016;
end
591876:begin
	ram_in<=32'd2016;
end
591877:begin
	ram_in<=32'd4064;
end
591878:begin
	ram_in<=32'd3680;
end
591879:begin
	ram_in<=32'd3696;
end
591880:begin
	ram_in<=32'd3696;
end
591881:begin
	ram_in<=32'd3696;
end
591882:begin
	ram_in<=32'd7920;
end
591883:begin
	ram_in<=32'd4080;
end
591884:begin
	ram_in<=32'd4088;
end
591885:begin
	ram_in<=32'd4088;
end
591886:begin
	ram_in<=32'd4088;
end
591887:begin
	ram_in<=32'd4088;
end
591888:begin
	ram_in<=32'd952;
end
591889:begin
	ram_in<=32'd56;
end
591890:begin
	ram_in<=32'd56;
end
591891:begin
	ram_in<=32'd56;
end
591892:begin
	ram_in<=32'd56;
end
591893:begin
	ram_in<=32'd56;
end
591894:begin
	ram_in<=32'd24;
end
591895:begin
	ram_in<=32'd56;
end
591896:begin
	ram_in<=32'd56;
end
591897:begin
	ram_in<=32'd56;
end
591898:begin
	ram_in<=32'd112;
end
591899:begin
	ram_in<=32'd1008;
end
591900:begin
	ram_in<=32'd2032;
end
591901:begin
	ram_in<=32'd1008;
end
591902:begin
	ram_in<=32'd992;
end
591903:begin
	ram_in<=32'd992;
end
592128:begin
	ram_in<=32'd112;
end
592129:begin
	ram_in<=32'd248;
end
592130:begin
	ram_in<=32'd504;
end
592131:begin
	ram_in<=32'd1020;
end
592132:begin
	ram_in<=32'd1016;
end
592133:begin
	ram_in<=32'd1976;
end
592134:begin
	ram_in<=32'd1816;
end
592135:begin
	ram_in<=32'd3896;
end
592136:begin
	ram_in<=32'd3632;
end
592137:begin
	ram_in<=32'd3632;
end
592138:begin
	ram_in<=32'd7216;
end
592139:begin
	ram_in<=32'd7200;
end
592140:begin
	ram_in<=32'd3640;
end
592141:begin
	ram_in<=32'd3640;
end
592142:begin
	ram_in<=32'd3896;
end
592143:begin
	ram_in<=32'd2032;
end
592144:begin
	ram_in<=32'd1008;
end
592145:begin
	ram_in<=32'd1008;
end
592146:begin
	ram_in<=32'd240;
end
592147:begin
	ram_in<=32'd112;
end
592148:begin
	ram_in<=32'd112;
end
592149:begin
	ram_in<=32'd224;
end
592150:begin
	ram_in<=32'd224;
end
592151:begin
	ram_in<=32'd448;
end
592152:begin
	ram_in<=32'd448;
end
592153:begin
	ram_in<=32'd448;
end
592154:begin
	ram_in<=32'd448;
end
592155:begin
	ram_in<=32'd448;
end
592156:begin
	ram_in<=32'd448;
end
592157:begin
	ram_in<=32'd448;
end
592158:begin
	ram_in<=32'd192;
end
592159:begin
	ram_in<=32'd192;
end
				endcase
			end
			else begin
				case({rlayer,rn,rin})
65536:begin
	ram_w<=32'd2147483651;
end
65537:begin
	ram_w<=32'd15;
end
65538:begin
	ram_w<=32'd5;
end
65539:begin
	ram_w<=32'd2147483671;
end
65540:begin
	ram_w<=32'd2147483662;
end
65541:begin
	ram_w<=32'd2147483652;
end
65542:begin
	ram_w<=32'd2147483671;
end
65543:begin
	ram_w<=32'd6;
end
65544:begin
	ram_w<=32'd13;
end
65545:begin
	ram_w<=32'd8;
end
65546:begin
	ram_w<=32'd2147483655;
end
65547:begin
	ram_w<=32'd21;
end
65548:begin
	ram_w<=32'd2147483649;
end
65549:begin
	ram_w<=32'd2147483662;
end
65550:begin
	ram_w<=32'd10;
end
65551:begin
	ram_w<=32'd2147483663;
end
65552:begin
	ram_w<=32'd2147483663;
end
65553:begin
	ram_w<=32'd7;
end
65554:begin
	ram_w<=32'd2;
end
65555:begin
	ram_w<=32'd2147483655;
end
65556:begin
	ram_w<=32'd1;
end
65557:begin
	ram_w<=32'd2147483652;
end
65558:begin
	ram_w<=32'd2147483662;
end
65559:begin
	ram_w<=32'd2147483652;
end
65560:begin
	ram_w<=32'd1;
end
65561:begin
	ram_w<=32'd9;
end
65562:begin
	ram_w<=32'd2147483659;
end
65563:begin
	ram_w<=32'd6;
end
65564:begin
	ram_w<=32'd5;
end
65565:begin
	ram_w<=32'd2147483657;
end
65566:begin
	ram_w<=32'd16;
end
65567:begin
	ram_w<=32'd13;
end
65568:begin
	ram_w<=32'd3;
end
65792:begin
	ram_w<=32'd2147483651;
end
65793:begin
	ram_w<=32'd2147483658;
end
65794:begin
	ram_w<=32'd5;
end
65795:begin
	ram_w<=32'd2;
end
65796:begin
	ram_w<=32'd2147483662;
end
65797:begin
	ram_w<=32'd3;
end
65798:begin
	ram_w<=32'd19;
end
65799:begin
	ram_w<=32'd2147483666;
end
65800:begin
	ram_w<=32'd2147483656;
end
65801:begin
	ram_w<=32'd2147483651;
end
65802:begin
	ram_w<=32'd0;
end
65803:begin
	ram_w<=32'd2147483650;
end
65804:begin
	ram_w<=32'd2147483657;
end
65805:begin
	ram_w<=32'd12;
end
65806:begin
	ram_w<=32'd6;
end
65807:begin
	ram_w<=32'd2147483658;
end
65808:begin
	ram_w<=32'd4;
end
65809:begin
	ram_w<=32'd2147483653;
end
65810:begin
	ram_w<=32'd2;
end
65811:begin
	ram_w<=32'd2147483656;
end
65812:begin
	ram_w<=32'd16;
end
65813:begin
	ram_w<=32'd2147483654;
end
65814:begin
	ram_w<=32'd2147483656;
end
65815:begin
	ram_w<=32'd2147483663;
end
65816:begin
	ram_w<=32'd11;
end
65817:begin
	ram_w<=32'd2147483659;
end
65818:begin
	ram_w<=32'd17;
end
65819:begin
	ram_w<=32'd2147483652;
end
65820:begin
	ram_w<=32'd5;
end
65821:begin
	ram_w<=32'd3;
end
65822:begin
	ram_w<=32'd9;
end
65823:begin
	ram_w<=32'd8;
end
65824:begin
	ram_w<=32'd2147483656;
end
66048:begin
	ram_w<=32'd2147483651;
end
66049:begin
	ram_w<=32'd5;
end
66050:begin
	ram_w<=32'd6;
end
66051:begin
	ram_w<=32'd2147483654;
end
66052:begin
	ram_w<=32'd2147483664;
end
66053:begin
	ram_w<=32'd5;
end
66054:begin
	ram_w<=32'd17;
end
66055:begin
	ram_w<=32'd2147483660;
end
66056:begin
	ram_w<=32'd3;
end
66057:begin
	ram_w<=32'd2147483656;
end
66058:begin
	ram_w<=32'd2147483664;
end
66059:begin
	ram_w<=32'd2147483670;
end
66060:begin
	ram_w<=32'd2147483665;
end
66061:begin
	ram_w<=32'd1;
end
66062:begin
	ram_w<=32'd2147483667;
end
66063:begin
	ram_w<=32'd2147483651;
end
66064:begin
	ram_w<=32'd2147483668;
end
66065:begin
	ram_w<=32'd1;
end
66066:begin
	ram_w<=32'd2147483664;
end
66067:begin
	ram_w<=32'd2147483652;
end
66068:begin
	ram_w<=32'd0;
end
66069:begin
	ram_w<=32'd1;
end
66070:begin
	ram_w<=32'd2147483657;
end
66071:begin
	ram_w<=32'd2147483655;
end
66072:begin
	ram_w<=32'd10;
end
66073:begin
	ram_w<=32'd0;
end
66074:begin
	ram_w<=32'd2147483649;
end
66075:begin
	ram_w<=32'd2147483666;
end
66076:begin
	ram_w<=32'd4;
end
66077:begin
	ram_w<=32'd2147483659;
end
66078:begin
	ram_w<=32'd7;
end
66079:begin
	ram_w<=32'd2147483654;
end
66080:begin
	ram_w<=32'd0;
end
66304:begin
	ram_w<=32'd0;
end
66305:begin
	ram_w<=32'd2;
end
66306:begin
	ram_w<=32'd13;
end
66307:begin
	ram_w<=32'd2147483652;
end
66308:begin
	ram_w<=32'd2147483655;
end
66309:begin
	ram_w<=32'd1;
end
66310:begin
	ram_w<=32'd2147483665;
end
66311:begin
	ram_w<=32'd2147483656;
end
66312:begin
	ram_w<=32'd9;
end
66313:begin
	ram_w<=32'd12;
end
66314:begin
	ram_w<=32'd2147483657;
end
66315:begin
	ram_w<=32'd2147483672;
end
66316:begin
	ram_w<=32'd1;
end
66317:begin
	ram_w<=32'd10;
end
66318:begin
	ram_w<=32'd2147483668;
end
66319:begin
	ram_w<=32'd2147483658;
end
66320:begin
	ram_w<=32'd2147483651;
end
66321:begin
	ram_w<=32'd19;
end
66322:begin
	ram_w<=32'd2147483656;
end
66323:begin
	ram_w<=32'd2147483670;
end
66324:begin
	ram_w<=32'd2147483655;
end
66325:begin
	ram_w<=32'd1;
end
66326:begin
	ram_w<=32'd2147483656;
end
66327:begin
	ram_w<=32'd22;
end
66328:begin
	ram_w<=32'd5;
end
66329:begin
	ram_w<=32'd2147483651;
end
66330:begin
	ram_w<=32'd2147483652;
end
66331:begin
	ram_w<=32'd2147483661;
end
66332:begin
	ram_w<=32'd2147483660;
end
66333:begin
	ram_w<=32'd2147483656;
end
66334:begin
	ram_w<=32'd8;
end
66335:begin
	ram_w<=32'd5;
end
66336:begin
	ram_w<=32'd2147483661;
end
66560:begin
	ram_w<=32'd6;
end
66561:begin
	ram_w<=32'd2147483649;
end
66562:begin
	ram_w<=32'd4;
end
66563:begin
	ram_w<=32'd2147483650;
end
66564:begin
	ram_w<=32'd3;
end
66565:begin
	ram_w<=32'd6;
end
66566:begin
	ram_w<=32'd8;
end
66567:begin
	ram_w<=32'd16;
end
66568:begin
	ram_w<=32'd2147483657;
end
66569:begin
	ram_w<=32'd2147483662;
end
66570:begin
	ram_w<=32'd2147483663;
end
66571:begin
	ram_w<=32'd2147483654;
end
66572:begin
	ram_w<=32'd2147483660;
end
66573:begin
	ram_w<=32'd7;
end
66574:begin
	ram_w<=32'd2147483649;
end
66575:begin
	ram_w<=32'd2147483652;
end
66576:begin
	ram_w<=32'd8;
end
66577:begin
	ram_w<=32'd7;
end
66578:begin
	ram_w<=32'd11;
end
66579:begin
	ram_w<=32'd2;
end
66580:begin
	ram_w<=32'd2147483652;
end
66581:begin
	ram_w<=32'd12;
end
66582:begin
	ram_w<=32'd2147483655;
end
66583:begin
	ram_w<=32'd8;
end
66584:begin
	ram_w<=32'd2147483651;
end
66585:begin
	ram_w<=32'd5;
end
66586:begin
	ram_w<=32'd2147483657;
end
66587:begin
	ram_w<=32'd2147483664;
end
66588:begin
	ram_w<=32'd0;
end
66589:begin
	ram_w<=32'd13;
end
66590:begin
	ram_w<=32'd0;
end
66591:begin
	ram_w<=32'd2147483665;
end
66592:begin
	ram_w<=32'd2147483651;
end
66816:begin
	ram_w<=32'd2147483653;
end
66817:begin
	ram_w<=32'd2147483655;
end
66818:begin
	ram_w<=32'd2147483651;
end
66819:begin
	ram_w<=32'd2;
end
66820:begin
	ram_w<=32'd5;
end
66821:begin
	ram_w<=32'd2147483662;
end
66822:begin
	ram_w<=32'd2147483651;
end
66823:begin
	ram_w<=32'd2147483658;
end
66824:begin
	ram_w<=32'd14;
end
66825:begin
	ram_w<=32'd2147483660;
end
66826:begin
	ram_w<=32'd2147483658;
end
66827:begin
	ram_w<=32'd6;
end
66828:begin
	ram_w<=32'd2147483658;
end
66829:begin
	ram_w<=32'd12;
end
66830:begin
	ram_w<=32'd2147483654;
end
66831:begin
	ram_w<=32'd7;
end
66832:begin
	ram_w<=32'd5;
end
66833:begin
	ram_w<=32'd2147483653;
end
66834:begin
	ram_w<=32'd7;
end
66835:begin
	ram_w<=32'd2147483652;
end
66836:begin
	ram_w<=32'd7;
end
66837:begin
	ram_w<=32'd5;
end
66838:begin
	ram_w<=32'd4;
end
66839:begin
	ram_w<=32'd22;
end
66840:begin
	ram_w<=32'd2147483660;
end
66841:begin
	ram_w<=32'd10;
end
66842:begin
	ram_w<=32'd2147483653;
end
66843:begin
	ram_w<=32'd2147483655;
end
66844:begin
	ram_w<=32'd7;
end
66845:begin
	ram_w<=32'd2147483664;
end
66846:begin
	ram_w<=32'd8;
end
66847:begin
	ram_w<=32'd2147483666;
end
66848:begin
	ram_w<=32'd5;
end
67072:begin
	ram_w<=32'd2147483656;
end
67073:begin
	ram_w<=32'd2147483667;
end
67074:begin
	ram_w<=32'd10;
end
67075:begin
	ram_w<=32'd2147483661;
end
67076:begin
	ram_w<=32'd2147483655;
end
67077:begin
	ram_w<=32'd2147483658;
end
67078:begin
	ram_w<=32'd17;
end
67079:begin
	ram_w<=32'd1;
end
67080:begin
	ram_w<=32'd2147483657;
end
67081:begin
	ram_w<=32'd2147483653;
end
67082:begin
	ram_w<=32'd2147483661;
end
67083:begin
	ram_w<=32'd2147483656;
end
67084:begin
	ram_w<=32'd0;
end
67085:begin
	ram_w<=32'd2;
end
67086:begin
	ram_w<=32'd9;
end
67087:begin
	ram_w<=32'd12;
end
67088:begin
	ram_w<=32'd8;
end
67089:begin
	ram_w<=32'd2147483659;
end
67090:begin
	ram_w<=32'd1;
end
67091:begin
	ram_w<=32'd2147483658;
end
67092:begin
	ram_w<=32'd2147483653;
end
67093:begin
	ram_w<=32'd5;
end
67094:begin
	ram_w<=32'd2147483651;
end
67095:begin
	ram_w<=32'd2147483652;
end
67096:begin
	ram_w<=32'd16;
end
67097:begin
	ram_w<=32'd2147483657;
end
67098:begin
	ram_w<=32'd2147483650;
end
67099:begin
	ram_w<=32'd2147483657;
end
67100:begin
	ram_w<=32'd2147483655;
end
67101:begin
	ram_w<=32'd2147483649;
end
67102:begin
	ram_w<=32'd2147483666;
end
67103:begin
	ram_w<=32'd2147483670;
end
67104:begin
	ram_w<=32'd2147483656;
end
67328:begin
	ram_w<=32'd2147483653;
end
67329:begin
	ram_w<=32'd6;
end
67330:begin
	ram_w<=32'd7;
end
67331:begin
	ram_w<=32'd2147483656;
end
67332:begin
	ram_w<=32'd17;
end
67333:begin
	ram_w<=32'd2147483670;
end
67334:begin
	ram_w<=32'd2147483659;
end
67335:begin
	ram_w<=32'd2147483670;
end
67336:begin
	ram_w<=32'd2147483667;
end
67337:begin
	ram_w<=32'd7;
end
67338:begin
	ram_w<=32'd2147483652;
end
67339:begin
	ram_w<=32'd1;
end
67340:begin
	ram_w<=32'd2147483658;
end
67341:begin
	ram_w<=32'd7;
end
67342:begin
	ram_w<=32'd14;
end
67343:begin
	ram_w<=32'd2147483660;
end
67344:begin
	ram_w<=32'd1;
end
67345:begin
	ram_w<=32'd0;
end
67346:begin
	ram_w<=32'd2147483651;
end
67347:begin
	ram_w<=32'd15;
end
67348:begin
	ram_w<=32'd2147483658;
end
67349:begin
	ram_w<=32'd2147483649;
end
67350:begin
	ram_w<=32'd2147483657;
end
67351:begin
	ram_w<=32'd14;
end
67352:begin
	ram_w<=32'd2147483650;
end
67353:begin
	ram_w<=32'd2147483656;
end
67354:begin
	ram_w<=32'd10;
end
67355:begin
	ram_w<=32'd1;
end
67356:begin
	ram_w<=32'd4;
end
67357:begin
	ram_w<=32'd1;
end
67358:begin
	ram_w<=32'd2147483654;
end
67359:begin
	ram_w<=32'd2147483653;
end
67360:begin
	ram_w<=32'd2147483652;
end
67584:begin
	ram_w<=32'd3;
end
67585:begin
	ram_w<=32'd9;
end
67586:begin
	ram_w<=32'd2147483656;
end
67587:begin
	ram_w<=32'd0;
end
67588:begin
	ram_w<=32'd2147483653;
end
67589:begin
	ram_w<=32'd2147483658;
end
67590:begin
	ram_w<=32'd1;
end
67591:begin
	ram_w<=32'd2147483650;
end
67592:begin
	ram_w<=32'd5;
end
67593:begin
	ram_w<=32'd17;
end
67594:begin
	ram_w<=32'd2147483649;
end
67595:begin
	ram_w<=32'd2147483657;
end
67596:begin
	ram_w<=32'd2147483667;
end
67597:begin
	ram_w<=32'd13;
end
67598:begin
	ram_w<=32'd2147483656;
end
67599:begin
	ram_w<=32'd2147483649;
end
67600:begin
	ram_w<=32'd2147483662;
end
67601:begin
	ram_w<=32'd12;
end
67602:begin
	ram_w<=32'd23;
end
67603:begin
	ram_w<=32'd2147483667;
end
67604:begin
	ram_w<=32'd2147483657;
end
67605:begin
	ram_w<=32'd2147483664;
end
67606:begin
	ram_w<=32'd2147483663;
end
67607:begin
	ram_w<=32'd2147483656;
end
67608:begin
	ram_w<=32'd6;
end
67609:begin
	ram_w<=32'd2147483661;
end
67610:begin
	ram_w<=32'd1;
end
67611:begin
	ram_w<=32'd11;
end
67612:begin
	ram_w<=32'd11;
end
67613:begin
	ram_w<=32'd2147483649;
end
67614:begin
	ram_w<=32'd11;
end
67615:begin
	ram_w<=32'd2;
end
67616:begin
	ram_w<=32'd2147483656;
end
67840:begin
	ram_w<=32'd2147483655;
end
67841:begin
	ram_w<=32'd1;
end
67842:begin
	ram_w<=32'd2147483654;
end
67843:begin
	ram_w<=32'd2147483650;
end
67844:begin
	ram_w<=32'd10;
end
67845:begin
	ram_w<=32'd17;
end
67846:begin
	ram_w<=32'd2147483652;
end
67847:begin
	ram_w<=32'd2147483650;
end
67848:begin
	ram_w<=32'd2147483655;
end
67849:begin
	ram_w<=32'd2147483654;
end
67850:begin
	ram_w<=32'd9;
end
67851:begin
	ram_w<=32'd7;
end
67852:begin
	ram_w<=32'd12;
end
67853:begin
	ram_w<=32'd1;
end
67854:begin
	ram_w<=32'd3;
end
67855:begin
	ram_w<=32'd6;
end
67856:begin
	ram_w<=32'd6;
end
67857:begin
	ram_w<=32'd8;
end
67858:begin
	ram_w<=32'd2147483649;
end
67859:begin
	ram_w<=32'd13;
end
67860:begin
	ram_w<=32'd2147483650;
end
67861:begin
	ram_w<=32'd3;
end
67862:begin
	ram_w<=32'd2147483656;
end
67863:begin
	ram_w<=32'd2147483659;
end
67864:begin
	ram_w<=32'd7;
end
67865:begin
	ram_w<=32'd9;
end
67866:begin
	ram_w<=32'd2147483660;
end
67867:begin
	ram_w<=32'd7;
end
67868:begin
	ram_w<=32'd18;
end
67869:begin
	ram_w<=32'd2147483650;
end
67870:begin
	ram_w<=32'd2147483651;
end
67871:begin
	ram_w<=32'd2147483660;
end
67872:begin
	ram_w<=32'd18;
end
68096:begin
	ram_w<=32'd2147483651;
end
68097:begin
	ram_w<=32'd2147483658;
end
68098:begin
	ram_w<=32'd2147483653;
end
68099:begin
	ram_w<=32'd8;
end
68100:begin
	ram_w<=32'd1;
end
68101:begin
	ram_w<=32'd2147483656;
end
68102:begin
	ram_w<=32'd2147483674;
end
68103:begin
	ram_w<=32'd2147483658;
end
68104:begin
	ram_w<=32'd2147483658;
end
68105:begin
	ram_w<=32'd1;
end
68106:begin
	ram_w<=32'd7;
end
68107:begin
	ram_w<=32'd15;
end
68108:begin
	ram_w<=32'd2147483655;
end
68109:begin
	ram_w<=32'd2147483671;
end
68110:begin
	ram_w<=32'd2147483654;
end
68111:begin
	ram_w<=32'd5;
end
68112:begin
	ram_w<=32'd2147483651;
end
68113:begin
	ram_w<=32'd10;
end
68114:begin
	ram_w<=32'd13;
end
68115:begin
	ram_w<=32'd2147483666;
end
68116:begin
	ram_w<=32'd2147483670;
end
68117:begin
	ram_w<=32'd3;
end
68118:begin
	ram_w<=32'd2147483666;
end
68119:begin
	ram_w<=32'd1;
end
68120:begin
	ram_w<=32'd3;
end
68121:begin
	ram_w<=32'd17;
end
68122:begin
	ram_w<=32'd4;
end
68123:begin
	ram_w<=32'd2147483650;
end
68124:begin
	ram_w<=32'd2147483663;
end
68125:begin
	ram_w<=32'd2147483657;
end
68126:begin
	ram_w<=32'd2147483664;
end
68127:begin
	ram_w<=32'd15;
end
68128:begin
	ram_w<=32'd2147483657;
end
68352:begin
	ram_w<=32'd2147483653;
end
68353:begin
	ram_w<=32'd2147483652;
end
68354:begin
	ram_w<=32'd2147483651;
end
68355:begin
	ram_w<=32'd2147483649;
end
68356:begin
	ram_w<=32'd2147483649;
end
68357:begin
	ram_w<=32'd2147483655;
end
68358:begin
	ram_w<=32'd11;
end
68359:begin
	ram_w<=32'd2147483653;
end
68360:begin
	ram_w<=32'd0;
end
68361:begin
	ram_w<=32'd17;
end
68362:begin
	ram_w<=32'd7;
end
68363:begin
	ram_w<=32'd2147483661;
end
68364:begin
	ram_w<=32'd15;
end
68365:begin
	ram_w<=32'd2147483656;
end
68366:begin
	ram_w<=32'd8;
end
68367:begin
	ram_w<=32'd0;
end
68368:begin
	ram_w<=32'd2147483655;
end
68369:begin
	ram_w<=32'd2147483653;
end
68370:begin
	ram_w<=32'd2147483650;
end
68371:begin
	ram_w<=32'd2147483649;
end
68372:begin
	ram_w<=32'd2147483667;
end
68373:begin
	ram_w<=32'd2147483654;
end
68374:begin
	ram_w<=32'd9;
end
68375:begin
	ram_w<=32'd2147483655;
end
68376:begin
	ram_w<=32'd7;
end
68377:begin
	ram_w<=32'd0;
end
68378:begin
	ram_w<=32'd4;
end
68379:begin
	ram_w<=32'd2147483667;
end
68380:begin
	ram_w<=32'd17;
end
68381:begin
	ram_w<=32'd2147483649;
end
68382:begin
	ram_w<=32'd8;
end
68383:begin
	ram_w<=32'd13;
end
68384:begin
	ram_w<=32'd2147483662;
end
68608:begin
	ram_w<=32'd0;
end
68609:begin
	ram_w<=32'd20;
end
68610:begin
	ram_w<=32'd14;
end
68611:begin
	ram_w<=32'd2;
end
68612:begin
	ram_w<=32'd2147483657;
end
68613:begin
	ram_w<=32'd19;
end
68614:begin
	ram_w<=32'd2147483654;
end
68615:begin
	ram_w<=32'd2147483666;
end
68616:begin
	ram_w<=32'd2147483665;
end
68617:begin
	ram_w<=32'd7;
end
68618:begin
	ram_w<=32'd2147483651;
end
68619:begin
	ram_w<=32'd0;
end
68620:begin
	ram_w<=32'd2147483653;
end
68621:begin
	ram_w<=32'd2147483662;
end
68622:begin
	ram_w<=32'd2147483661;
end
68623:begin
	ram_w<=32'd2147483656;
end
68624:begin
	ram_w<=32'd2147483661;
end
68625:begin
	ram_w<=32'd2147483653;
end
68626:begin
	ram_w<=32'd6;
end
68627:begin
	ram_w<=32'd2147483656;
end
68628:begin
	ram_w<=32'd1;
end
68629:begin
	ram_w<=32'd2;
end
68630:begin
	ram_w<=32'd9;
end
68631:begin
	ram_w<=32'd0;
end
68632:begin
	ram_w<=32'd2147483654;
end
68633:begin
	ram_w<=32'd3;
end
68634:begin
	ram_w<=32'd2147483657;
end
68635:begin
	ram_w<=32'd6;
end
68636:begin
	ram_w<=32'd7;
end
68637:begin
	ram_w<=32'd2147483653;
end
68638:begin
	ram_w<=32'd2147483650;
end
68639:begin
	ram_w<=32'd2147483662;
end
68640:begin
	ram_w<=32'd13;
end
68864:begin
	ram_w<=32'd2147483649;
end
68865:begin
	ram_w<=32'd22;
end
68866:begin
	ram_w<=32'd1;
end
68867:begin
	ram_w<=32'd13;
end
68868:begin
	ram_w<=32'd1;
end
68869:begin
	ram_w<=32'd6;
end
68870:begin
	ram_w<=32'd19;
end
68871:begin
	ram_w<=32'd2;
end
68872:begin
	ram_w<=32'd2147483662;
end
68873:begin
	ram_w<=32'd2147483664;
end
68874:begin
	ram_w<=32'd2147483654;
end
68875:begin
	ram_w<=32'd2147483672;
end
68876:begin
	ram_w<=32'd2147483659;
end
68877:begin
	ram_w<=32'd2147483654;
end
68878:begin
	ram_w<=32'd2147483653;
end
68879:begin
	ram_w<=32'd2147483651;
end
68880:begin
	ram_w<=32'd0;
end
68881:begin
	ram_w<=32'd0;
end
68882:begin
	ram_w<=32'd2147483651;
end
68883:begin
	ram_w<=32'd6;
end
68884:begin
	ram_w<=32'd2147483652;
end
68885:begin
	ram_w<=32'd4;
end
68886:begin
	ram_w<=32'd16;
end
68887:begin
	ram_w<=32'd5;
end
68888:begin
	ram_w<=32'd2;
end
68889:begin
	ram_w<=32'd2147483655;
end
68890:begin
	ram_w<=32'd4;
end
68891:begin
	ram_w<=32'd0;
end
68892:begin
	ram_w<=32'd2147483655;
end
68893:begin
	ram_w<=32'd5;
end
68894:begin
	ram_w<=32'd2147483657;
end
68895:begin
	ram_w<=32'd2147483659;
end
68896:begin
	ram_w<=32'd6;
end
69120:begin
	ram_w<=32'd4;
end
69121:begin
	ram_w<=32'd17;
end
69122:begin
	ram_w<=32'd4;
end
69123:begin
	ram_w<=32'd14;
end
69124:begin
	ram_w<=32'd2147483651;
end
69125:begin
	ram_w<=32'd17;
end
69126:begin
	ram_w<=32'd2147483661;
end
69127:begin
	ram_w<=32'd0;
end
69128:begin
	ram_w<=32'd1;
end
69129:begin
	ram_w<=32'd3;
end
69130:begin
	ram_w<=32'd3;
end
69131:begin
	ram_w<=32'd9;
end
69132:begin
	ram_w<=32'd3;
end
69133:begin
	ram_w<=32'd14;
end
69134:begin
	ram_w<=32'd3;
end
69135:begin
	ram_w<=32'd8;
end
69136:begin
	ram_w<=32'd12;
end
69137:begin
	ram_w<=32'd3;
end
69138:begin
	ram_w<=32'd20;
end
69139:begin
	ram_w<=32'd2147483650;
end
69140:begin
	ram_w<=32'd0;
end
69141:begin
	ram_w<=32'd7;
end
69142:begin
	ram_w<=32'd13;
end
69143:begin
	ram_w<=32'd16;
end
69144:begin
	ram_w<=32'd2147483649;
end
69145:begin
	ram_w<=32'd6;
end
69146:begin
	ram_w<=32'd2147483658;
end
69147:begin
	ram_w<=32'd2147483654;
end
69148:begin
	ram_w<=32'd11;
end
69149:begin
	ram_w<=32'd2147483656;
end
69150:begin
	ram_w<=32'd2147483667;
end
69151:begin
	ram_w<=32'd2147483653;
end
69152:begin
	ram_w<=32'd3;
end
69376:begin
	ram_w<=32'd0;
end
69377:begin
	ram_w<=32'd2147483659;
end
69378:begin
	ram_w<=32'd2147483649;
end
69379:begin
	ram_w<=32'd5;
end
69380:begin
	ram_w<=32'd3;
end
69381:begin
	ram_w<=32'd11;
end
69382:begin
	ram_w<=32'd9;
end
69383:begin
	ram_w<=32'd2147483668;
end
69384:begin
	ram_w<=32'd2147483665;
end
69385:begin
	ram_w<=32'd2147483660;
end
69386:begin
	ram_w<=32'd18;
end
69387:begin
	ram_w<=32'd2147483664;
end
69388:begin
	ram_w<=32'd3;
end
69389:begin
	ram_w<=32'd2147483655;
end
69390:begin
	ram_w<=32'd2147483651;
end
69391:begin
	ram_w<=32'd8;
end
69392:begin
	ram_w<=32'd11;
end
69393:begin
	ram_w<=32'd2147483653;
end
69394:begin
	ram_w<=32'd7;
end
69395:begin
	ram_w<=32'd0;
end
69396:begin
	ram_w<=32'd11;
end
69397:begin
	ram_w<=32'd1;
end
69398:begin
	ram_w<=32'd2147483665;
end
69399:begin
	ram_w<=32'd1;
end
69400:begin
	ram_w<=32'd6;
end
69401:begin
	ram_w<=32'd2147483657;
end
69402:begin
	ram_w<=32'd3;
end
69403:begin
	ram_w<=32'd2147483661;
end
69404:begin
	ram_w<=32'd0;
end
69405:begin
	ram_w<=32'd2147483659;
end
69406:begin
	ram_w<=32'd2147483657;
end
69407:begin
	ram_w<=32'd2147483653;
end
69408:begin
	ram_w<=32'd4;
end
69632:begin
	ram_w<=32'd2147483655;
end
69633:begin
	ram_w<=32'd2147483653;
end
69634:begin
	ram_w<=32'd4;
end
69635:begin
	ram_w<=32'd2147483653;
end
69636:begin
	ram_w<=32'd2147483652;
end
69637:begin
	ram_w<=32'd2147483651;
end
69638:begin
	ram_w<=32'd2147483651;
end
69639:begin
	ram_w<=32'd2147483661;
end
69640:begin
	ram_w<=32'd2147483673;
end
69641:begin
	ram_w<=32'd1;
end
69642:begin
	ram_w<=32'd2147483658;
end
69643:begin
	ram_w<=32'd2147483655;
end
69644:begin
	ram_w<=32'd2147483666;
end
69645:begin
	ram_w<=32'd9;
end
69646:begin
	ram_w<=32'd2147483655;
end
69647:begin
	ram_w<=32'd2;
end
69648:begin
	ram_w<=32'd7;
end
69649:begin
	ram_w<=32'd0;
end
69650:begin
	ram_w<=32'd2147483657;
end
69651:begin
	ram_w<=32'd8;
end
69652:begin
	ram_w<=32'd2147483660;
end
69653:begin
	ram_w<=32'd1;
end
69654:begin
	ram_w<=32'd17;
end
69655:begin
	ram_w<=32'd1;
end
69656:begin
	ram_w<=32'd3;
end
69657:begin
	ram_w<=32'd2;
end
69658:begin
	ram_w<=32'd0;
end
69659:begin
	ram_w<=32'd7;
end
69660:begin
	ram_w<=32'd2147483654;
end
69661:begin
	ram_w<=32'd4;
end
69662:begin
	ram_w<=32'd3;
end
69663:begin
	ram_w<=32'd2147483658;
end
69664:begin
	ram_w<=32'd8;
end
69888:begin
	ram_w<=32'd0;
end
69889:begin
	ram_w<=32'd2147483652;
end
69890:begin
	ram_w<=32'd12;
end
69891:begin
	ram_w<=32'd2147483653;
end
69892:begin
	ram_w<=32'd9;
end
69893:begin
	ram_w<=32'd13;
end
69894:begin
	ram_w<=32'd0;
end
69895:begin
	ram_w<=32'd9;
end
69896:begin
	ram_w<=32'd0;
end
69897:begin
	ram_w<=32'd5;
end
69898:begin
	ram_w<=32'd2147483656;
end
69899:begin
	ram_w<=32'd2147483649;
end
69900:begin
	ram_w<=32'd7;
end
69901:begin
	ram_w<=32'd2147483651;
end
69902:begin
	ram_w<=32'd0;
end
69903:begin
	ram_w<=32'd4;
end
69904:begin
	ram_w<=32'd5;
end
69905:begin
	ram_w<=32'd2147483651;
end
69906:begin
	ram_w<=32'd2147483653;
end
69907:begin
	ram_w<=32'd4;
end
69908:begin
	ram_w<=32'd3;
end
69909:begin
	ram_w<=32'd0;
end
69910:begin
	ram_w<=32'd2147483652;
end
69911:begin
	ram_w<=32'd2147483652;
end
69912:begin
	ram_w<=32'd2147483662;
end
69913:begin
	ram_w<=32'd2147483651;
end
69914:begin
	ram_w<=32'd2147483659;
end
69915:begin
	ram_w<=32'd2147483653;
end
69916:begin
	ram_w<=32'd0;
end
69917:begin
	ram_w<=32'd2147483653;
end
69918:begin
	ram_w<=32'd4;
end
69919:begin
	ram_w<=32'd2147483654;
end
69920:begin
	ram_w<=32'd7;
end
70144:begin
	ram_w<=32'd2147483652;
end
70145:begin
	ram_w<=32'd2147483665;
end
70146:begin
	ram_w<=32'd2147483660;
end
70147:begin
	ram_w<=32'd14;
end
70148:begin
	ram_w<=32'd5;
end
70149:begin
	ram_w<=32'd2147483671;
end
70150:begin
	ram_w<=32'd2147483654;
end
70151:begin
	ram_w<=32'd2147483663;
end
70152:begin
	ram_w<=32'd3;
end
70153:begin
	ram_w<=32'd4;
end
70154:begin
	ram_w<=32'd2147483651;
end
70155:begin
	ram_w<=32'd2147483652;
end
70156:begin
	ram_w<=32'd14;
end
70157:begin
	ram_w<=32'd2147483654;
end
70158:begin
	ram_w<=32'd3;
end
70159:begin
	ram_w<=32'd3;
end
70160:begin
	ram_w<=32'd4;
end
70161:begin
	ram_w<=32'd2147483653;
end
70162:begin
	ram_w<=32'd2147483660;
end
70163:begin
	ram_w<=32'd2147483653;
end
70164:begin
	ram_w<=32'd2147483656;
end
70165:begin
	ram_w<=32'd2147483654;
end
70166:begin
	ram_w<=32'd2147483649;
end
70167:begin
	ram_w<=32'd16;
end
70168:begin
	ram_w<=32'd4;
end
70169:begin
	ram_w<=32'd2147483652;
end
70170:begin
	ram_w<=32'd2147483652;
end
70171:begin
	ram_w<=32'd2147483651;
end
70172:begin
	ram_w<=32'd3;
end
70173:begin
	ram_w<=32'd4;
end
70174:begin
	ram_w<=32'd8;
end
70175:begin
	ram_w<=32'd2147483651;
end
70176:begin
	ram_w<=32'd7;
end
70400:begin
	ram_w<=32'd2147483653;
end
70401:begin
	ram_w<=32'd5;
end
70402:begin
	ram_w<=32'd2147483660;
end
70403:begin
	ram_w<=32'd5;
end
70404:begin
	ram_w<=32'd2147483651;
end
70405:begin
	ram_w<=32'd2147483667;
end
70406:begin
	ram_w<=32'd6;
end
70407:begin
	ram_w<=32'd3;
end
70408:begin
	ram_w<=32'd2147483662;
end
70409:begin
	ram_w<=32'd17;
end
70410:begin
	ram_w<=32'd2147483653;
end
70411:begin
	ram_w<=32'd1;
end
70412:begin
	ram_w<=32'd2147483663;
end
70413:begin
	ram_w<=32'd17;
end
70414:begin
	ram_w<=32'd2147483652;
end
70415:begin
	ram_w<=32'd2147483652;
end
70416:begin
	ram_w<=32'd2147483655;
end
70417:begin
	ram_w<=32'd2147483664;
end
70418:begin
	ram_w<=32'd2147483659;
end
70419:begin
	ram_w<=32'd2147483655;
end
70420:begin
	ram_w<=32'd2147483661;
end
70421:begin
	ram_w<=32'd2147483655;
end
70422:begin
	ram_w<=32'd2147483654;
end
70423:begin
	ram_w<=32'd7;
end
70424:begin
	ram_w<=32'd2147483651;
end
70425:begin
	ram_w<=32'd2147483666;
end
70426:begin
	ram_w<=32'd2147483651;
end
70427:begin
	ram_w<=32'd11;
end
70428:begin
	ram_w<=32'd13;
end
70429:begin
	ram_w<=32'd2147483653;
end
70430:begin
	ram_w<=32'd17;
end
70431:begin
	ram_w<=32'd2147483652;
end
70432:begin
	ram_w<=32'd2147483657;
end
70656:begin
	ram_w<=32'd2147483652;
end
70657:begin
	ram_w<=32'd7;
end
70658:begin
	ram_w<=32'd2147483656;
end
70659:begin
	ram_w<=32'd2147483660;
end
70660:begin
	ram_w<=32'd2147483656;
end
70661:begin
	ram_w<=32'd2147483649;
end
70662:begin
	ram_w<=32'd2147483652;
end
70663:begin
	ram_w<=32'd4;
end
70664:begin
	ram_w<=32'd4;
end
70665:begin
	ram_w<=32'd4;
end
70666:begin
	ram_w<=32'd7;
end
70667:begin
	ram_w<=32'd12;
end
70668:begin
	ram_w<=32'd2147483662;
end
70669:begin
	ram_w<=32'd11;
end
70670:begin
	ram_w<=32'd4;
end
70671:begin
	ram_w<=32'd2147483652;
end
70672:begin
	ram_w<=32'd6;
end
70673:begin
	ram_w<=32'd11;
end
70674:begin
	ram_w<=32'd17;
end
70675:begin
	ram_w<=32'd2147483661;
end
70676:begin
	ram_w<=32'd2147483659;
end
70677:begin
	ram_w<=32'd13;
end
70678:begin
	ram_w<=32'd6;
end
70679:begin
	ram_w<=32'd15;
end
70680:begin
	ram_w<=32'd2147483651;
end
70681:begin
	ram_w<=32'd2147483649;
end
70682:begin
	ram_w<=32'd2147483656;
end
70683:begin
	ram_w<=32'd1;
end
70684:begin
	ram_w<=32'd3;
end
70685:begin
	ram_w<=32'd1;
end
70686:begin
	ram_w<=32'd2147483650;
end
70687:begin
	ram_w<=32'd2147483650;
end
70688:begin
	ram_w<=32'd2147483651;
end
70912:begin
	ram_w<=32'd2147483650;
end
70913:begin
	ram_w<=32'd9;
end
70914:begin
	ram_w<=32'd2147483656;
end
70915:begin
	ram_w<=32'd7;
end
70916:begin
	ram_w<=32'd17;
end
70917:begin
	ram_w<=32'd2147483658;
end
70918:begin
	ram_w<=32'd2147483654;
end
70919:begin
	ram_w<=32'd0;
end
70920:begin
	ram_w<=32'd2147483656;
end
70921:begin
	ram_w<=32'd2147483660;
end
70922:begin
	ram_w<=32'd2147483654;
end
70923:begin
	ram_w<=32'd2147483651;
end
70924:begin
	ram_w<=32'd2147483651;
end
70925:begin
	ram_w<=32'd2147483650;
end
70926:begin
	ram_w<=32'd8;
end
70927:begin
	ram_w<=32'd2147483654;
end
70928:begin
	ram_w<=32'd2147483657;
end
70929:begin
	ram_w<=32'd2147483667;
end
70930:begin
	ram_w<=32'd2147483653;
end
70931:begin
	ram_w<=32'd11;
end
70932:begin
	ram_w<=32'd2147483653;
end
70933:begin
	ram_w<=32'd1;
end
70934:begin
	ram_w<=32'd2147483653;
end
70935:begin
	ram_w<=32'd2147483659;
end
70936:begin
	ram_w<=32'd4;
end
70937:begin
	ram_w<=32'd7;
end
70938:begin
	ram_w<=32'd2;
end
70939:begin
	ram_w<=32'd2147483660;
end
70940:begin
	ram_w<=32'd10;
end
70941:begin
	ram_w<=32'd2147483653;
end
70942:begin
	ram_w<=32'd2147483663;
end
70943:begin
	ram_w<=32'd1;
end
70944:begin
	ram_w<=32'd5;
end
71168:begin
	ram_w<=32'd2147483650;
end
71169:begin
	ram_w<=32'd2147483662;
end
71170:begin
	ram_w<=32'd2147483657;
end
71171:begin
	ram_w<=32'd2;
end
71172:begin
	ram_w<=32'd2147483668;
end
71173:begin
	ram_w<=32'd2147483669;
end
71174:begin
	ram_w<=32'd2147483649;
end
71175:begin
	ram_w<=32'd2147483654;
end
71176:begin
	ram_w<=32'd2147483670;
end
71177:begin
	ram_w<=32'd0;
end
71178:begin
	ram_w<=32'd2147483650;
end
71179:begin
	ram_w<=32'd2147483664;
end
71180:begin
	ram_w<=32'd5;
end
71181:begin
	ram_w<=32'd2;
end
71182:begin
	ram_w<=32'd2147483654;
end
71183:begin
	ram_w<=32'd17;
end
71184:begin
	ram_w<=32'd5;
end
71185:begin
	ram_w<=32'd6;
end
71186:begin
	ram_w<=32'd2147483651;
end
71187:begin
	ram_w<=32'd2147483652;
end
71188:begin
	ram_w<=32'd3;
end
71189:begin
	ram_w<=32'd2147483658;
end
71190:begin
	ram_w<=32'd1;
end
71191:begin
	ram_w<=32'd1;
end
71192:begin
	ram_w<=32'd2147483665;
end
71193:begin
	ram_w<=32'd2147483650;
end
71194:begin
	ram_w<=32'd2147483662;
end
71195:begin
	ram_w<=32'd2147483653;
end
71196:begin
	ram_w<=32'd2147483649;
end
71197:begin
	ram_w<=32'd0;
end
71198:begin
	ram_w<=32'd19;
end
71199:begin
	ram_w<=32'd6;
end
71200:begin
	ram_w<=32'd2147483660;
end
71424:begin
	ram_w<=32'd2147483651;
end
71425:begin
	ram_w<=32'd2147483654;
end
71426:begin
	ram_w<=32'd11;
end
71427:begin
	ram_w<=32'd5;
end
71428:begin
	ram_w<=32'd16;
end
71429:begin
	ram_w<=32'd2147483667;
end
71430:begin
	ram_w<=32'd13;
end
71431:begin
	ram_w<=32'd3;
end
71432:begin
	ram_w<=32'd4;
end
71433:begin
	ram_w<=32'd2147483658;
end
71434:begin
	ram_w<=32'd2147483656;
end
71435:begin
	ram_w<=32'd2147483650;
end
71436:begin
	ram_w<=32'd2147483663;
end
71437:begin
	ram_w<=32'd12;
end
71438:begin
	ram_w<=32'd8;
end
71439:begin
	ram_w<=32'd12;
end
71440:begin
	ram_w<=32'd2147483651;
end
71441:begin
	ram_w<=32'd2147483649;
end
71442:begin
	ram_w<=32'd2147483669;
end
71443:begin
	ram_w<=32'd2147483658;
end
71444:begin
	ram_w<=32'd2147483663;
end
71445:begin
	ram_w<=32'd10;
end
71446:begin
	ram_w<=32'd2147483659;
end
71447:begin
	ram_w<=32'd2;
end
71448:begin
	ram_w<=32'd5;
end
71449:begin
	ram_w<=32'd2147483656;
end
71450:begin
	ram_w<=32'd9;
end
71451:begin
	ram_w<=32'd2147483653;
end
71452:begin
	ram_w<=32'd0;
end
71453:begin
	ram_w<=32'd2147483655;
end
71454:begin
	ram_w<=32'd2147483665;
end
71455:begin
	ram_w<=32'd0;
end
71456:begin
	ram_w<=32'd2147483653;
end
71680:begin
	ram_w<=32'd4;
end
71681:begin
	ram_w<=32'd12;
end
71682:begin
	ram_w<=32'd2147483665;
end
71683:begin
	ram_w<=32'd2147483655;
end
71684:begin
	ram_w<=32'd2147483651;
end
71685:begin
	ram_w<=32'd2147483670;
end
71686:begin
	ram_w<=32'd2147483664;
end
71687:begin
	ram_w<=32'd2147483657;
end
71688:begin
	ram_w<=32'd3;
end
71689:begin
	ram_w<=32'd2147483668;
end
71690:begin
	ram_w<=32'd2147483653;
end
71691:begin
	ram_w<=32'd3;
end
71692:begin
	ram_w<=32'd15;
end
71693:begin
	ram_w<=32'd2;
end
71694:begin
	ram_w<=32'd2147483654;
end
71695:begin
	ram_w<=32'd5;
end
71696:begin
	ram_w<=32'd13;
end
71697:begin
	ram_w<=32'd2147483649;
end
71698:begin
	ram_w<=32'd2147483656;
end
71699:begin
	ram_w<=32'd1;
end
71700:begin
	ram_w<=32'd11;
end
71701:begin
	ram_w<=32'd2147483658;
end
71702:begin
	ram_w<=32'd4;
end
71703:begin
	ram_w<=32'd2147483654;
end
71704:begin
	ram_w<=32'd1;
end
71705:begin
	ram_w<=32'd9;
end
71706:begin
	ram_w<=32'd1;
end
71707:begin
	ram_w<=32'd2147483666;
end
71708:begin
	ram_w<=32'd1;
end
71709:begin
	ram_w<=32'd2147483667;
end
71710:begin
	ram_w<=32'd0;
end
71711:begin
	ram_w<=32'd6;
end
71712:begin
	ram_w<=32'd20;
end
71936:begin
	ram_w<=32'd7;
end
71937:begin
	ram_w<=32'd2147483666;
end
71938:begin
	ram_w<=32'd2147483673;
end
71939:begin
	ram_w<=32'd2147483650;
end
71940:begin
	ram_w<=32'd8;
end
71941:begin
	ram_w<=32'd2147483650;
end
71942:begin
	ram_w<=32'd13;
end
71943:begin
	ram_w<=32'd2147483649;
end
71944:begin
	ram_w<=32'd15;
end
71945:begin
	ram_w<=32'd4;
end
71946:begin
	ram_w<=32'd5;
end
71947:begin
	ram_w<=32'd10;
end
71948:begin
	ram_w<=32'd11;
end
71949:begin
	ram_w<=32'd2147483650;
end
71950:begin
	ram_w<=32'd8;
end
71951:begin
	ram_w<=32'd6;
end
71952:begin
	ram_w<=32'd3;
end
71953:begin
	ram_w<=32'd2147483657;
end
71954:begin
	ram_w<=32'd2147483658;
end
71955:begin
	ram_w<=32'd11;
end
71956:begin
	ram_w<=32'd2147483659;
end
71957:begin
	ram_w<=32'd0;
end
71958:begin
	ram_w<=32'd0;
end
71959:begin
	ram_w<=32'd2147483649;
end
71960:begin
	ram_w<=32'd0;
end
71961:begin
	ram_w<=32'd4;
end
71962:begin
	ram_w<=32'd7;
end
71963:begin
	ram_w<=32'd15;
end
71964:begin
	ram_w<=32'd13;
end
71965:begin
	ram_w<=32'd3;
end
71966:begin
	ram_w<=32'd10;
end
71967:begin
	ram_w<=32'd2147483667;
end
71968:begin
	ram_w<=32'd2147483655;
end
72192:begin
	ram_w<=32'd1;
end
72193:begin
	ram_w<=32'd2147483656;
end
72194:begin
	ram_w<=32'd2147483651;
end
72195:begin
	ram_w<=32'd21;
end
72196:begin
	ram_w<=32'd5;
end
72197:begin
	ram_w<=32'd2147483649;
end
72198:begin
	ram_w<=32'd5;
end
72199:begin
	ram_w<=32'd2147483661;
end
72200:begin
	ram_w<=32'd2147483649;
end
72201:begin
	ram_w<=32'd2147483653;
end
72202:begin
	ram_w<=32'd2147483649;
end
72203:begin
	ram_w<=32'd3;
end
72204:begin
	ram_w<=32'd10;
end
72205:begin
	ram_w<=32'd4;
end
72206:begin
	ram_w<=32'd6;
end
72207:begin
	ram_w<=32'd2147483651;
end
72208:begin
	ram_w<=32'd2147483649;
end
72209:begin
	ram_w<=32'd8;
end
72210:begin
	ram_w<=32'd12;
end
72211:begin
	ram_w<=32'd1;
end
72212:begin
	ram_w<=32'd2147483649;
end
72213:begin
	ram_w<=32'd2147483654;
end
72214:begin
	ram_w<=32'd17;
end
72215:begin
	ram_w<=32'd2147483649;
end
72216:begin
	ram_w<=32'd2147483656;
end
72217:begin
	ram_w<=32'd13;
end
72218:begin
	ram_w<=32'd12;
end
72219:begin
	ram_w<=32'd2147483649;
end
72220:begin
	ram_w<=32'd0;
end
72221:begin
	ram_w<=32'd4;
end
72222:begin
	ram_w<=32'd2147483661;
end
72223:begin
	ram_w<=32'd2147483654;
end
72224:begin
	ram_w<=32'd15;
end
72448:begin
	ram_w<=32'd2147483651;
end
72449:begin
	ram_w<=32'd8;
end
72450:begin
	ram_w<=32'd1;
end
72451:begin
	ram_w<=32'd2147483664;
end
72452:begin
	ram_w<=32'd2147483649;
end
72453:begin
	ram_w<=32'd5;
end
72454:begin
	ram_w<=32'd2147483663;
end
72455:begin
	ram_w<=32'd2147483658;
end
72456:begin
	ram_w<=32'd2147483662;
end
72457:begin
	ram_w<=32'd2147483652;
end
72458:begin
	ram_w<=32'd2147483657;
end
72459:begin
	ram_w<=32'd2147483656;
end
72460:begin
	ram_w<=32'd2147483661;
end
72461:begin
	ram_w<=32'd5;
end
72462:begin
	ram_w<=32'd7;
end
72463:begin
	ram_w<=32'd3;
end
72464:begin
	ram_w<=32'd9;
end
72465:begin
	ram_w<=32'd4;
end
72466:begin
	ram_w<=32'd2147483668;
end
72467:begin
	ram_w<=32'd2147483669;
end
72468:begin
	ram_w<=32'd2147483662;
end
72469:begin
	ram_w<=32'd2147483662;
end
72470:begin
	ram_w<=32'd3;
end
72471:begin
	ram_w<=32'd2147483668;
end
72472:begin
	ram_w<=32'd8;
end
72473:begin
	ram_w<=32'd2147483667;
end
72474:begin
	ram_w<=32'd5;
end
72475:begin
	ram_w<=32'd2147483668;
end
72476:begin
	ram_w<=32'd2147483659;
end
72477:begin
	ram_w<=32'd2147483659;
end
72478:begin
	ram_w<=32'd0;
end
72479:begin
	ram_w<=32'd2147483658;
end
72480:begin
	ram_w<=32'd12;
end
72704:begin
	ram_w<=32'd2147483652;
end
72705:begin
	ram_w<=32'd13;
end
72706:begin
	ram_w<=32'd4;
end
72707:begin
	ram_w<=32'd2147483654;
end
72708:begin
	ram_w<=32'd2147483651;
end
72709:begin
	ram_w<=32'd8;
end
72710:begin
	ram_w<=32'd2147483649;
end
72711:begin
	ram_w<=32'd4;
end
72712:begin
	ram_w<=32'd2147483650;
end
72713:begin
	ram_w<=32'd2147483649;
end
72714:begin
	ram_w<=32'd2;
end
72715:begin
	ram_w<=32'd2147483657;
end
72716:begin
	ram_w<=32'd2147483650;
end
72717:begin
	ram_w<=32'd2147483649;
end
72718:begin
	ram_w<=32'd2147483655;
end
72719:begin
	ram_w<=32'd4;
end
72720:begin
	ram_w<=32'd2147483652;
end
72721:begin
	ram_w<=32'd2147483649;
end
72722:begin
	ram_w<=32'd15;
end
72723:begin
	ram_w<=32'd2;
end
72724:begin
	ram_w<=32'd0;
end
72725:begin
	ram_w<=32'd2147483656;
end
72726:begin
	ram_w<=32'd11;
end
72727:begin
	ram_w<=32'd5;
end
72728:begin
	ram_w<=32'd2147483657;
end
72729:begin
	ram_w<=32'd13;
end
72730:begin
	ram_w<=32'd3;
end
72731:begin
	ram_w<=32'd2147483656;
end
72732:begin
	ram_w<=32'd2147483652;
end
72733:begin
	ram_w<=32'd10;
end
72734:begin
	ram_w<=32'd7;
end
72735:begin
	ram_w<=32'd2147483661;
end
72736:begin
	ram_w<=32'd2147483650;
end
72960:begin
	ram_w<=32'd1;
end
72961:begin
	ram_w<=32'd2147483662;
end
72962:begin
	ram_w<=32'd13;
end
72963:begin
	ram_w<=32'd7;
end
72964:begin
	ram_w<=32'd9;
end
72965:begin
	ram_w<=32'd1;
end
72966:begin
	ram_w<=32'd2147483652;
end
72967:begin
	ram_w<=32'd2147483651;
end
72968:begin
	ram_w<=32'd2147483650;
end
72969:begin
	ram_w<=32'd10;
end
72970:begin
	ram_w<=32'd9;
end
72971:begin
	ram_w<=32'd7;
end
72972:begin
	ram_w<=32'd6;
end
72973:begin
	ram_w<=32'd2147483661;
end
72974:begin
	ram_w<=32'd2147483653;
end
72975:begin
	ram_w<=32'd2147483653;
end
72976:begin
	ram_w<=32'd7;
end
72977:begin
	ram_w<=32'd2147483658;
end
72978:begin
	ram_w<=32'd2147483663;
end
72979:begin
	ram_w<=32'd2147483659;
end
72980:begin
	ram_w<=32'd2147483668;
end
72981:begin
	ram_w<=32'd15;
end
72982:begin
	ram_w<=32'd2;
end
72983:begin
	ram_w<=32'd2147483649;
end
72984:begin
	ram_w<=32'd2147483654;
end
72985:begin
	ram_w<=32'd2147483655;
end
72986:begin
	ram_w<=32'd2147483660;
end
72987:begin
	ram_w<=32'd2147483669;
end
72988:begin
	ram_w<=32'd2147483651;
end
72989:begin
	ram_w<=32'd2147483663;
end
72990:begin
	ram_w<=32'd2147483661;
end
72991:begin
	ram_w<=32'd1;
end
72992:begin
	ram_w<=32'd5;
end
131072:begin
	ram_w<=32'd2147483661;
end
131073:begin
	ram_w<=32'd2147483659;
end
131074:begin
	ram_w<=32'd8;
end
131075:begin
	ram_w<=32'd10;
end
131076:begin
	ram_w<=32'd17;
end
131077:begin
	ram_w<=32'd2147483657;
end
131078:begin
	ram_w<=32'd9;
end
131079:begin
	ram_w<=32'd2147483649;
end
131080:begin
	ram_w<=32'd6;
end
131081:begin
	ram_w<=32'd2147483649;
end
131082:begin
	ram_w<=32'd0;
end
131083:begin
	ram_w<=32'd2147483663;
end
131084:begin
	ram_w<=32'd2147483654;
end
131085:begin
	ram_w<=32'd7;
end
131086:begin
	ram_w<=32'd2147483663;
end
131087:begin
	ram_w<=32'd9;
end
131088:begin
	ram_w<=32'd2147483654;
end
131089:begin
	ram_w<=32'd2147483660;
end
131090:begin
	ram_w<=32'd2147483659;
end
131091:begin
	ram_w<=32'd2147483651;
end
131092:begin
	ram_w<=32'd4;
end
131093:begin
	ram_w<=32'd6;
end
131094:begin
	ram_w<=32'd4;
end
131095:begin
	ram_w<=32'd2147483651;
end
131096:begin
	ram_w<=32'd2147483652;
end
131097:begin
	ram_w<=32'd2147483666;
end
131098:begin
	ram_w<=32'd3;
end
131099:begin
	ram_w<=32'd2147483654;
end
131100:begin
	ram_w<=32'd2147483649;
end
131101:begin
	ram_w<=32'd12;
end
131102:begin
	ram_w<=32'd2;
end
131328:begin
	ram_w<=32'd9;
end
131329:begin
	ram_w<=32'd3;
end
131330:begin
	ram_w<=32'd1;
end
131331:begin
	ram_w<=32'd3;
end
131332:begin
	ram_w<=32'd2147483655;
end
131333:begin
	ram_w<=32'd8;
end
131334:begin
	ram_w<=32'd2147483654;
end
131335:begin
	ram_w<=32'd2147483658;
end
131336:begin
	ram_w<=32'd2147483649;
end
131337:begin
	ram_w<=32'd0;
end
131338:begin
	ram_w<=32'd2147483660;
end
131339:begin
	ram_w<=32'd1;
end
131340:begin
	ram_w<=32'd2147483649;
end
131341:begin
	ram_w<=32'd0;
end
131342:begin
	ram_w<=32'd2147483660;
end
131343:begin
	ram_w<=32'd15;
end
131344:begin
	ram_w<=32'd0;
end
131345:begin
	ram_w<=32'd2147483651;
end
131346:begin
	ram_w<=32'd2147483661;
end
131347:begin
	ram_w<=32'd7;
end
131348:begin
	ram_w<=32'd12;
end
131349:begin
	ram_w<=32'd2147483650;
end
131350:begin
	ram_w<=32'd4;
end
131351:begin
	ram_w<=32'd10;
end
131352:begin
	ram_w<=32'd13;
end
131353:begin
	ram_w<=32'd8;
end
131354:begin
	ram_w<=32'd4;
end
131355:begin
	ram_w<=32'd6;
end
131356:begin
	ram_w<=32'd2;
end
131357:begin
	ram_w<=32'd2147483650;
end
131358:begin
	ram_w<=32'd1;
end
131584:begin
	ram_w<=32'd2147483651;
end
131585:begin
	ram_w<=32'd2147483650;
end
131586:begin
	ram_w<=32'd2147483657;
end
131587:begin
	ram_w<=32'd11;
end
131588:begin
	ram_w<=32'd2147483649;
end
131589:begin
	ram_w<=32'd2147483658;
end
131590:begin
	ram_w<=32'd8;
end
131591:begin
	ram_w<=32'd10;
end
131592:begin
	ram_w<=32'd8;
end
131593:begin
	ram_w<=32'd2147483654;
end
131594:begin
	ram_w<=32'd2;
end
131595:begin
	ram_w<=32'd2147483650;
end
131596:begin
	ram_w<=32'd8;
end
131597:begin
	ram_w<=32'd2147483654;
end
131598:begin
	ram_w<=32'd3;
end
131599:begin
	ram_w<=32'd1;
end
131600:begin
	ram_w<=32'd2147483659;
end
131601:begin
	ram_w<=32'd2147483655;
end
131602:begin
	ram_w<=32'd0;
end
131603:begin
	ram_w<=32'd2147483650;
end
131604:begin
	ram_w<=32'd3;
end
131605:begin
	ram_w<=32'd5;
end
131606:begin
	ram_w<=32'd14;
end
131607:begin
	ram_w<=32'd2147483654;
end
131608:begin
	ram_w<=32'd2147483650;
end
131609:begin
	ram_w<=32'd2147483662;
end
131610:begin
	ram_w<=32'd2;
end
131611:begin
	ram_w<=32'd3;
end
131612:begin
	ram_w<=32'd2147483649;
end
131613:begin
	ram_w<=32'd12;
end
131614:begin
	ram_w<=32'd2147483653;
end
131840:begin
	ram_w<=32'd1;
end
131841:begin
	ram_w<=32'd2147483652;
end
131842:begin
	ram_w<=32'd1;
end
131843:begin
	ram_w<=32'd2147483656;
end
131844:begin
	ram_w<=32'd2147483656;
end
131845:begin
	ram_w<=32'd3;
end
131846:begin
	ram_w<=32'd2147483658;
end
131847:begin
	ram_w<=32'd2147483658;
end
131848:begin
	ram_w<=32'd3;
end
131849:begin
	ram_w<=32'd5;
end
131850:begin
	ram_w<=32'd8;
end
131851:begin
	ram_w<=32'd2147483649;
end
131852:begin
	ram_w<=32'd4;
end
131853:begin
	ram_w<=32'd7;
end
131854:begin
	ram_w<=32'd2147483658;
end
131855:begin
	ram_w<=32'd2147483658;
end
131856:begin
	ram_w<=32'd7;
end
131857:begin
	ram_w<=32'd2147483656;
end
131858:begin
	ram_w<=32'd4;
end
131859:begin
	ram_w<=32'd9;
end
131860:begin
	ram_w<=32'd2147483658;
end
131861:begin
	ram_w<=32'd15;
end
131862:begin
	ram_w<=32'd5;
end
131863:begin
	ram_w<=32'd2147483656;
end
131864:begin
	ram_w<=32'd16;
end
131865:begin
	ram_w<=32'd1;
end
131866:begin
	ram_w<=32'd2147483649;
end
131867:begin
	ram_w<=32'd2;
end
131868:begin
	ram_w<=32'd2147483665;
end
131869:begin
	ram_w<=32'd9;
end
131870:begin
	ram_w<=32'd3;
end
132096:begin
	ram_w<=32'd2147483653;
end
132097:begin
	ram_w<=32'd2147483663;
end
132098:begin
	ram_w<=32'd2147483660;
end
132099:begin
	ram_w<=32'd2147483650;
end
132100:begin
	ram_w<=32'd2147483658;
end
132101:begin
	ram_w<=32'd2147483658;
end
132102:begin
	ram_w<=32'd14;
end
132103:begin
	ram_w<=32'd2147483660;
end
132104:begin
	ram_w<=32'd12;
end
132105:begin
	ram_w<=32'd2147483652;
end
132106:begin
	ram_w<=32'd2147483653;
end
132107:begin
	ram_w<=32'd2147483653;
end
132108:begin
	ram_w<=32'd5;
end
132109:begin
	ram_w<=32'd2147483654;
end
132110:begin
	ram_w<=32'd2147483662;
end
132111:begin
	ram_w<=32'd2147483650;
end
132112:begin
	ram_w<=32'd6;
end
132113:begin
	ram_w<=32'd18;
end
132114:begin
	ram_w<=32'd11;
end
132115:begin
	ram_w<=32'd12;
end
132116:begin
	ram_w<=32'd3;
end
132117:begin
	ram_w<=32'd15;
end
132118:begin
	ram_w<=32'd2147483653;
end
132119:begin
	ram_w<=32'd2147483649;
end
132120:begin
	ram_w<=32'd2147483654;
end
132121:begin
	ram_w<=32'd7;
end
132122:begin
	ram_w<=32'd2147483650;
end
132123:begin
	ram_w<=32'd15;
end
132124:begin
	ram_w<=32'd2147483656;
end
132125:begin
	ram_w<=32'd2147483650;
end
132126:begin
	ram_w<=32'd2147483662;
end
132352:begin
	ram_w<=32'd2147483651;
end
132353:begin
	ram_w<=32'd2147483654;
end
132354:begin
	ram_w<=32'd2147483652;
end
132355:begin
	ram_w<=32'd2147483655;
end
132356:begin
	ram_w<=32'd17;
end
132357:begin
	ram_w<=32'd2;
end
132358:begin
	ram_w<=32'd3;
end
132359:begin
	ram_w<=32'd2147483658;
end
132360:begin
	ram_w<=32'd2147483655;
end
132361:begin
	ram_w<=32'd0;
end
132362:begin
	ram_w<=32'd4;
end
132363:begin
	ram_w<=32'd2147483655;
end
132364:begin
	ram_w<=32'd7;
end
132365:begin
	ram_w<=32'd9;
end
132366:begin
	ram_w<=32'd2147483668;
end
132367:begin
	ram_w<=32'd3;
end
132368:begin
	ram_w<=32'd2147483655;
end
132369:begin
	ram_w<=32'd8;
end
132370:begin
	ram_w<=32'd0;
end
132371:begin
	ram_w<=32'd2147483660;
end
132372:begin
	ram_w<=32'd2147483651;
end
132373:begin
	ram_w<=32'd3;
end
132374:begin
	ram_w<=32'd2;
end
132375:begin
	ram_w<=32'd7;
end
132376:begin
	ram_w<=32'd5;
end
132377:begin
	ram_w<=32'd2147483651;
end
132378:begin
	ram_w<=32'd0;
end
132379:begin
	ram_w<=32'd4;
end
132380:begin
	ram_w<=32'd2147483652;
end
132381:begin
	ram_w<=32'd2147483650;
end
132382:begin
	ram_w<=32'd2147483649;
end
132608:begin
	ram_w<=32'd10;
end
132609:begin
	ram_w<=32'd2147483671;
end
132610:begin
	ram_w<=32'd5;
end
132611:begin
	ram_w<=32'd2147483671;
end
132612:begin
	ram_w<=32'd8;
end
132613:begin
	ram_w<=32'd2147483659;
end
132614:begin
	ram_w<=32'd15;
end
132615:begin
	ram_w<=32'd2147483659;
end
132616:begin
	ram_w<=32'd6;
end
132617:begin
	ram_w<=32'd2147483659;
end
132618:begin
	ram_w<=32'd5;
end
132619:begin
	ram_w<=32'd2147483649;
end
132620:begin
	ram_w<=32'd2147483657;
end
132621:begin
	ram_w<=32'd11;
end
132622:begin
	ram_w<=32'd2147483672;
end
132623:begin
	ram_w<=32'd7;
end
132624:begin
	ram_w<=32'd2147483665;
end
132625:begin
	ram_w<=32'd5;
end
132626:begin
	ram_w<=32'd2147483663;
end
132627:begin
	ram_w<=32'd2147483650;
end
132628:begin
	ram_w<=32'd3;
end
132629:begin
	ram_w<=32'd9;
end
132630:begin
	ram_w<=32'd9;
end
132631:begin
	ram_w<=32'd2147483660;
end
132632:begin
	ram_w<=32'd2147483657;
end
132633:begin
	ram_w<=32'd2147483655;
end
132634:begin
	ram_w<=32'd2;
end
132635:begin
	ram_w<=32'd2147483657;
end
132636:begin
	ram_w<=32'd5;
end
132637:begin
	ram_w<=32'd16;
end
132638:begin
	ram_w<=32'd2147483658;
end
132864:begin
	ram_w<=32'd6;
end
132865:begin
	ram_w<=32'd2147483659;
end
132866:begin
	ram_w<=32'd2147483654;
end
132867:begin
	ram_w<=32'd15;
end
132868:begin
	ram_w<=32'd14;
end
132869:begin
	ram_w<=32'd2;
end
132870:begin
	ram_w<=32'd2147483654;
end
132871:begin
	ram_w<=32'd2147483661;
end
132872:begin
	ram_w<=32'd8;
end
132873:begin
	ram_w<=32'd4;
end
132874:begin
	ram_w<=32'd2147483657;
end
132875:begin
	ram_w<=32'd2147483666;
end
132876:begin
	ram_w<=32'd1;
end
132877:begin
	ram_w<=32'd3;
end
132878:begin
	ram_w<=32'd2147483649;
end
132879:begin
	ram_w<=32'd9;
end
132880:begin
	ram_w<=32'd7;
end
132881:begin
	ram_w<=32'd8;
end
132882:begin
	ram_w<=32'd4;
end
132883:begin
	ram_w<=32'd12;
end
132884:begin
	ram_w<=32'd8;
end
132885:begin
	ram_w<=32'd2147483653;
end
132886:begin
	ram_w<=32'd2147483664;
end
132887:begin
	ram_w<=32'd16;
end
132888:begin
	ram_w<=32'd6;
end
132889:begin
	ram_w<=32'd2147483655;
end
132890:begin
	ram_w<=32'd2;
end
132891:begin
	ram_w<=32'd9;
end
132892:begin
	ram_w<=32'd1;
end
132893:begin
	ram_w<=32'd3;
end
132894:begin
	ram_w<=32'd14;
end
133120:begin
	ram_w<=32'd2147483649;
end
133121:begin
	ram_w<=32'd2147483653;
end
133122:begin
	ram_w<=32'd2147483654;
end
133123:begin
	ram_w<=32'd9;
end
133124:begin
	ram_w<=32'd2147483652;
end
133125:begin
	ram_w<=32'd2147483657;
end
133126:begin
	ram_w<=32'd9;
end
133127:begin
	ram_w<=32'd6;
end
133128:begin
	ram_w<=32'd2147483661;
end
133129:begin
	ram_w<=32'd2147483675;
end
133130:begin
	ram_w<=32'd2147483656;
end
133131:begin
	ram_w<=32'd2147483658;
end
133132:begin
	ram_w<=32'd2;
end
133133:begin
	ram_w<=32'd7;
end
133134:begin
	ram_w<=32'd2147483652;
end
133135:begin
	ram_w<=32'd5;
end
133136:begin
	ram_w<=32'd0;
end
133137:begin
	ram_w<=32'd2147483650;
end
133138:begin
	ram_w<=32'd4;
end
133139:begin
	ram_w<=32'd2147483654;
end
133140:begin
	ram_w<=32'd9;
end
133141:begin
	ram_w<=32'd6;
end
133142:begin
	ram_w<=32'd2147483659;
end
133143:begin
	ram_w<=32'd6;
end
133144:begin
	ram_w<=32'd2147483656;
end
133145:begin
	ram_w<=32'd2147483663;
end
133146:begin
	ram_w<=32'd5;
end
133147:begin
	ram_w<=32'd10;
end
133148:begin
	ram_w<=32'd18;
end
133149:begin
	ram_w<=32'd3;
end
133150:begin
	ram_w<=32'd2147483655;
end
133376:begin
	ram_w<=32'd6;
end
133377:begin
	ram_w<=32'd2147483661;
end
133378:begin
	ram_w<=32'd5;
end
133379:begin
	ram_w<=32'd2147483654;
end
133380:begin
	ram_w<=32'd1;
end
133381:begin
	ram_w<=32'd2147483656;
end
133382:begin
	ram_w<=32'd7;
end
133383:begin
	ram_w<=32'd2147483651;
end
133384:begin
	ram_w<=32'd11;
end
133385:begin
	ram_w<=32'd2147483653;
end
133386:begin
	ram_w<=32'd2147483654;
end
133387:begin
	ram_w<=32'd12;
end
133388:begin
	ram_w<=32'd2147483649;
end
133389:begin
	ram_w<=32'd2147483655;
end
133390:begin
	ram_w<=32'd2147483652;
end
133391:begin
	ram_w<=32'd1;
end
133392:begin
	ram_w<=32'd0;
end
133393:begin
	ram_w<=32'd2;
end
133394:begin
	ram_w<=32'd8;
end
133395:begin
	ram_w<=32'd7;
end
133396:begin
	ram_w<=32'd9;
end
133397:begin
	ram_w<=32'd11;
end
133398:begin
	ram_w<=32'd18;
end
133399:begin
	ram_w<=32'd2147483649;
end
133400:begin
	ram_w<=32'd2147483652;
end
133401:begin
	ram_w<=32'd4;
end
133402:begin
	ram_w<=32'd5;
end
133403:begin
	ram_w<=32'd8;
end
133404:begin
	ram_w<=32'd2147483649;
end
133405:begin
	ram_w<=32'd2147483658;
end
133406:begin
	ram_w<=32'd7;
end
				endcase
			end
			rf<=1;
			state<=IDLE;
		end
		endcase
	end
end

endmodule

