module connect#(
parameter maxl=5,
parameter sizein=32,
parameter sizew=8,
parameter sizeout=40
)
(
input clk,
input rst,
input start,

output reg[7:0] rlayer,//the layer to be read
output reg[7:0] rn,//the neuron to be read
output reg[7:0] rin,//the input of a neuron
output reg rmode,//0: read input, 1: read weight/bias
output reg rs,//start
input[sizein-1:0] ram_in,
input[sizew-1:0] ram_w,
input rf,//finished

output reg[7:0] result,
output reg finished,
output [31:0] debug,
output [31:0] debug1,
output [sizeout-1:0] prob0,
output [sizeout-1:0] prob1,
output [sizeout-1:0] prob2,
output [sizeout-1:0] prob3,
output [sizeout-1:0] out0,
output [sizeout-1:0] out1,
output [sizeout-1:0] out2,
output [sizeout-1:0] out3,
output [sizeout-1:0] out4,
output [sizeout-1:0] out5,
output [sizeout-1:0] out6,
output [sizeout-1:0] out7,
output [sizeout-1:0] out8,
output [sizeout-1:0] out9
);

reg[sizein-1:0] in[31:0];
reg[sizew-1:0] w[1:0][29:0][31:0];
reg[sizew-1:0] b[1:0][29:0];
wire[sizeout-1:0] out[29:0];
reg [sizeout-1:0] outtemp[29:0];
reg relu;

assign prob0=w[0][1][2];
assign prob1=b[0][2];
assign prob2=w[1][2][3];
assign prob3=b[1][4];

assign out0=out[0];
assign out1=out[1];
assign out2=out[2];
assign out3=out[3];
assign out4=out[4];
assign out5=out[5];
assign out6=out[6];
assign out7=out[7];
assign out8=out[8];
assign out9=out[9];

neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_0(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][0][0],w[0][0][1],w[0][0][2],w[0][0][3],w[0][0][4],w[0][0][5],w[0][0][6],w[0][0][7],w[0][0][8],w[0][0][9],w[0][0][10],w[0][0][11],w[0][0][12],w[0][0][13],w[0][0][14],w[0][0][15],w[0][0][16],w[0][0][17],w[0][0][18],w[0][0][19],w[0][0][20],w[0][0][21],w[0][0][22],w[0][0][23],w[0][0][24],w[0][0][25],w[0][0][26],w[0][0][27],w[0][0][28],w[0][0][29],w[0][0][30],w[0][0][31],b[0][0],out[0]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_1(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][1][0],w[0][1][1],w[0][1][2],w[0][1][3],w[0][1][4],w[0][1][5],w[0][1][6],w[0][1][7],w[0][1][8],w[0][1][9],w[0][1][10],w[0][1][11],w[0][1][12],w[0][1][13],w[0][1][14],w[0][1][15],w[0][1][16],w[0][1][17],w[0][1][18],w[0][1][19],w[0][1][20],w[0][1][21],w[0][1][22],w[0][1][23],w[0][1][24],w[0][1][25],w[0][1][26],w[0][1][27],w[0][1][28],w[0][1][29],w[0][1][30],w[0][1][31],b[0][1],out[1]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_2(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][2][0],w[0][2][1],w[0][2][2],w[0][2][3],w[0][2][4],w[0][2][5],w[0][2][6],w[0][2][7],w[0][2][8],w[0][2][9],w[0][2][10],w[0][2][11],w[0][2][12],w[0][2][13],w[0][2][14],w[0][2][15],w[0][2][16],w[0][2][17],w[0][2][18],w[0][2][19],w[0][2][20],w[0][2][21],w[0][2][22],w[0][2][23],w[0][2][24],w[0][2][25],w[0][2][26],w[0][2][27],w[0][2][28],w[0][2][29],w[0][2][30],w[0][2][31],b[0][2],out[2]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_3(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][3][0],w[0][3][1],w[0][3][2],w[0][3][3],w[0][3][4],w[0][3][5],w[0][3][6],w[0][3][7],w[0][3][8],w[0][3][9],w[0][3][10],w[0][3][11],w[0][3][12],w[0][3][13],w[0][3][14],w[0][3][15],w[0][3][16],w[0][3][17],w[0][3][18],w[0][3][19],w[0][3][20],w[0][3][21],w[0][3][22],w[0][3][23],w[0][3][24],w[0][3][25],w[0][3][26],w[0][3][27],w[0][3][28],w[0][3][29],w[0][3][30],w[0][3][31],b[0][3],out[3]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_4(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][4][0],w[0][4][1],w[0][4][2],w[0][4][3],w[0][4][4],w[0][4][5],w[0][4][6],w[0][4][7],w[0][4][8],w[0][4][9],w[0][4][10],w[0][4][11],w[0][4][12],w[0][4][13],w[0][4][14],w[0][4][15],w[0][4][16],w[0][4][17],w[0][4][18],w[0][4][19],w[0][4][20],w[0][4][21],w[0][4][22],w[0][4][23],w[0][4][24],w[0][4][25],w[0][4][26],w[0][4][27],w[0][4][28],w[0][4][29],w[0][4][30],w[0][4][31],b[0][4],out[4]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_5(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][5][0],w[0][5][1],w[0][5][2],w[0][5][3],w[0][5][4],w[0][5][5],w[0][5][6],w[0][5][7],w[0][5][8],w[0][5][9],w[0][5][10],w[0][5][11],w[0][5][12],w[0][5][13],w[0][5][14],w[0][5][15],w[0][5][16],w[0][5][17],w[0][5][18],w[0][5][19],w[0][5][20],w[0][5][21],w[0][5][22],w[0][5][23],w[0][5][24],w[0][5][25],w[0][5][26],w[0][5][27],w[0][5][28],w[0][5][29],w[0][5][30],w[0][5][31],b[0][5],out[5]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_6(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][6][0],w[0][6][1],w[0][6][2],w[0][6][3],w[0][6][4],w[0][6][5],w[0][6][6],w[0][6][7],w[0][6][8],w[0][6][9],w[0][6][10],w[0][6][11],w[0][6][12],w[0][6][13],w[0][6][14],w[0][6][15],w[0][6][16],w[0][6][17],w[0][6][18],w[0][6][19],w[0][6][20],w[0][6][21],w[0][6][22],w[0][6][23],w[0][6][24],w[0][6][25],w[0][6][26],w[0][6][27],w[0][6][28],w[0][6][29],w[0][6][30],w[0][6][31],b[0][6],out[6]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_7(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][7][0],w[0][7][1],w[0][7][2],w[0][7][3],w[0][7][4],w[0][7][5],w[0][7][6],w[0][7][7],w[0][7][8],w[0][7][9],w[0][7][10],w[0][7][11],w[0][7][12],w[0][7][13],w[0][7][14],w[0][7][15],w[0][7][16],w[0][7][17],w[0][7][18],w[0][7][19],w[0][7][20],w[0][7][21],w[0][7][22],w[0][7][23],w[0][7][24],w[0][7][25],w[0][7][26],w[0][7][27],w[0][7][28],w[0][7][29],w[0][7][30],w[0][7][31],b[0][7],out[7]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_8(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][8][0],w[0][8][1],w[0][8][2],w[0][8][3],w[0][8][4],w[0][8][5],w[0][8][6],w[0][8][7],w[0][8][8],w[0][8][9],w[0][8][10],w[0][8][11],w[0][8][12],w[0][8][13],w[0][8][14],w[0][8][15],w[0][8][16],w[0][8][17],w[0][8][18],w[0][8][19],w[0][8][20],w[0][8][21],w[0][8][22],w[0][8][23],w[0][8][24],w[0][8][25],w[0][8][26],w[0][8][27],w[0][8][28],w[0][8][29],w[0][8][30],w[0][8][31],b[0][8],out[8]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_9(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][9][0],w[0][9][1],w[0][9][2],w[0][9][3],w[0][9][4],w[0][9][5],w[0][9][6],w[0][9][7],w[0][9][8],w[0][9][9],w[0][9][10],w[0][9][11],w[0][9][12],w[0][9][13],w[0][9][14],w[0][9][15],w[0][9][16],w[0][9][17],w[0][9][18],w[0][9][19],w[0][9][20],w[0][9][21],w[0][9][22],w[0][9][23],w[0][9][24],w[0][9][25],w[0][9][26],w[0][9][27],w[0][9][28],w[0][9][29],w[0][9][30],w[0][9][31],b[0][9],out[9]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_10(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][10][0],w[0][10][1],w[0][10][2],w[0][10][3],w[0][10][4],w[0][10][5],w[0][10][6],w[0][10][7],w[0][10][8],w[0][10][9],w[0][10][10],w[0][10][11],w[0][10][12],w[0][10][13],w[0][10][14],w[0][10][15],w[0][10][16],w[0][10][17],w[0][10][18],w[0][10][19],w[0][10][20],w[0][10][21],w[0][10][22],w[0][10][23],w[0][10][24],w[0][10][25],w[0][10][26],w[0][10][27],w[0][10][28],w[0][10][29],w[0][10][30],w[0][10][31],b[0][10],out[10]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_11(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][11][0],w[0][11][1],w[0][11][2],w[0][11][3],w[0][11][4],w[0][11][5],w[0][11][6],w[0][11][7],w[0][11][8],w[0][11][9],w[0][11][10],w[0][11][11],w[0][11][12],w[0][11][13],w[0][11][14],w[0][11][15],w[0][11][16],w[0][11][17],w[0][11][18],w[0][11][19],w[0][11][20],w[0][11][21],w[0][11][22],w[0][11][23],w[0][11][24],w[0][11][25],w[0][11][26],w[0][11][27],w[0][11][28],w[0][11][29],w[0][11][30],w[0][11][31],b[0][11],out[11]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_12(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][12][0],w[0][12][1],w[0][12][2],w[0][12][3],w[0][12][4],w[0][12][5],w[0][12][6],w[0][12][7],w[0][12][8],w[0][12][9],w[0][12][10],w[0][12][11],w[0][12][12],w[0][12][13],w[0][12][14],w[0][12][15],w[0][12][16],w[0][12][17],w[0][12][18],w[0][12][19],w[0][12][20],w[0][12][21],w[0][12][22],w[0][12][23],w[0][12][24],w[0][12][25],w[0][12][26],w[0][12][27],w[0][12][28],w[0][12][29],w[0][12][30],w[0][12][31],b[0][12],out[12]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_13(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][13][0],w[0][13][1],w[0][13][2],w[0][13][3],w[0][13][4],w[0][13][5],w[0][13][6],w[0][13][7],w[0][13][8],w[0][13][9],w[0][13][10],w[0][13][11],w[0][13][12],w[0][13][13],w[0][13][14],w[0][13][15],w[0][13][16],w[0][13][17],w[0][13][18],w[0][13][19],w[0][13][20],w[0][13][21],w[0][13][22],w[0][13][23],w[0][13][24],w[0][13][25],w[0][13][26],w[0][13][27],w[0][13][28],w[0][13][29],w[0][13][30],w[0][13][31],b[0][13],out[13]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_14(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][14][0],w[0][14][1],w[0][14][2],w[0][14][3],w[0][14][4],w[0][14][5],w[0][14][6],w[0][14][7],w[0][14][8],w[0][14][9],w[0][14][10],w[0][14][11],w[0][14][12],w[0][14][13],w[0][14][14],w[0][14][15],w[0][14][16],w[0][14][17],w[0][14][18],w[0][14][19],w[0][14][20],w[0][14][21],w[0][14][22],w[0][14][23],w[0][14][24],w[0][14][25],w[0][14][26],w[0][14][27],w[0][14][28],w[0][14][29],w[0][14][30],w[0][14][31],b[0][14],out[14]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_15(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][15][0],w[0][15][1],w[0][15][2],w[0][15][3],w[0][15][4],w[0][15][5],w[0][15][6],w[0][15][7],w[0][15][8],w[0][15][9],w[0][15][10],w[0][15][11],w[0][15][12],w[0][15][13],w[0][15][14],w[0][15][15],w[0][15][16],w[0][15][17],w[0][15][18],w[0][15][19],w[0][15][20],w[0][15][21],w[0][15][22],w[0][15][23],w[0][15][24],w[0][15][25],w[0][15][26],w[0][15][27],w[0][15][28],w[0][15][29],w[0][15][30],w[0][15][31],b[0][15],out[15]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_16(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][16][0],w[0][16][1],w[0][16][2],w[0][16][3],w[0][16][4],w[0][16][5],w[0][16][6],w[0][16][7],w[0][16][8],w[0][16][9],w[0][16][10],w[0][16][11],w[0][16][12],w[0][16][13],w[0][16][14],w[0][16][15],w[0][16][16],w[0][16][17],w[0][16][18],w[0][16][19],w[0][16][20],w[0][16][21],w[0][16][22],w[0][16][23],w[0][16][24],w[0][16][25],w[0][16][26],w[0][16][27],w[0][16][28],w[0][16][29],w[0][16][30],w[0][16][31],b[0][16],out[16]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_17(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][17][0],w[0][17][1],w[0][17][2],w[0][17][3],w[0][17][4],w[0][17][5],w[0][17][6],w[0][17][7],w[0][17][8],w[0][17][9],w[0][17][10],w[0][17][11],w[0][17][12],w[0][17][13],w[0][17][14],w[0][17][15],w[0][17][16],w[0][17][17],w[0][17][18],w[0][17][19],w[0][17][20],w[0][17][21],w[0][17][22],w[0][17][23],w[0][17][24],w[0][17][25],w[0][17][26],w[0][17][27],w[0][17][28],w[0][17][29],w[0][17][30],w[0][17][31],b[0][17],out[17]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_18(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][18][0],w[0][18][1],w[0][18][2],w[0][18][3],w[0][18][4],w[0][18][5],w[0][18][6],w[0][18][7],w[0][18][8],w[0][18][9],w[0][18][10],w[0][18][11],w[0][18][12],w[0][18][13],w[0][18][14],w[0][18][15],w[0][18][16],w[0][18][17],w[0][18][18],w[0][18][19],w[0][18][20],w[0][18][21],w[0][18][22],w[0][18][23],w[0][18][24],w[0][18][25],w[0][18][26],w[0][18][27],w[0][18][28],w[0][18][29],w[0][18][30],w[0][18][31],b[0][18],out[18]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_19(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][19][0],w[0][19][1],w[0][19][2],w[0][19][3],w[0][19][4],w[0][19][5],w[0][19][6],w[0][19][7],w[0][19][8],w[0][19][9],w[0][19][10],w[0][19][11],w[0][19][12],w[0][19][13],w[0][19][14],w[0][19][15],w[0][19][16],w[0][19][17],w[0][19][18],w[0][19][19],w[0][19][20],w[0][19][21],w[0][19][22],w[0][19][23],w[0][19][24],w[0][19][25],w[0][19][26],w[0][19][27],w[0][19][28],w[0][19][29],w[0][19][30],w[0][19][31],b[0][19],out[19]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_20(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][20][0],w[0][20][1],w[0][20][2],w[0][20][3],w[0][20][4],w[0][20][5],w[0][20][6],w[0][20][7],w[0][20][8],w[0][20][9],w[0][20][10],w[0][20][11],w[0][20][12],w[0][20][13],w[0][20][14],w[0][20][15],w[0][20][16],w[0][20][17],w[0][20][18],w[0][20][19],w[0][20][20],w[0][20][21],w[0][20][22],w[0][20][23],w[0][20][24],w[0][20][25],w[0][20][26],w[0][20][27],w[0][20][28],w[0][20][29],w[0][20][30],w[0][20][31],b[0][20],out[20]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_21(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][21][0],w[0][21][1],w[0][21][2],w[0][21][3],w[0][21][4],w[0][21][5],w[0][21][6],w[0][21][7],w[0][21][8],w[0][21][9],w[0][21][10],w[0][21][11],w[0][21][12],w[0][21][13],w[0][21][14],w[0][21][15],w[0][21][16],w[0][21][17],w[0][21][18],w[0][21][19],w[0][21][20],w[0][21][21],w[0][21][22],w[0][21][23],w[0][21][24],w[0][21][25],w[0][21][26],w[0][21][27],w[0][21][28],w[0][21][29],w[0][21][30],w[0][21][31],b[0][21],out[21]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_22(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][22][0],w[0][22][1],w[0][22][2],w[0][22][3],w[0][22][4],w[0][22][5],w[0][22][6],w[0][22][7],w[0][22][8],w[0][22][9],w[0][22][10],w[0][22][11],w[0][22][12],w[0][22][13],w[0][22][14],w[0][22][15],w[0][22][16],w[0][22][17],w[0][22][18],w[0][22][19],w[0][22][20],w[0][22][21],w[0][22][22],w[0][22][23],w[0][22][24],w[0][22][25],w[0][22][26],w[0][22][27],w[0][22][28],w[0][22][29],w[0][22][30],w[0][22][31],b[0][22],out[22]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_23(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][23][0],w[0][23][1],w[0][23][2],w[0][23][3],w[0][23][4],w[0][23][5],w[0][23][6],w[0][23][7],w[0][23][8],w[0][23][9],w[0][23][10],w[0][23][11],w[0][23][12],w[0][23][13],w[0][23][14],w[0][23][15],w[0][23][16],w[0][23][17],w[0][23][18],w[0][23][19],w[0][23][20],w[0][23][21],w[0][23][22],w[0][23][23],w[0][23][24],w[0][23][25],w[0][23][26],w[0][23][27],w[0][23][28],w[0][23][29],w[0][23][30],w[0][23][31],b[0][23],out[23]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_24(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][24][0],w[0][24][1],w[0][24][2],w[0][24][3],w[0][24][4],w[0][24][5],w[0][24][6],w[0][24][7],w[0][24][8],w[0][24][9],w[0][24][10],w[0][24][11],w[0][24][12],w[0][24][13],w[0][24][14],w[0][24][15],w[0][24][16],w[0][24][17],w[0][24][18],w[0][24][19],w[0][24][20],w[0][24][21],w[0][24][22],w[0][24][23],w[0][24][24],w[0][24][25],w[0][24][26],w[0][24][27],w[0][24][28],w[0][24][29],w[0][24][30],w[0][24][31],b[0][24],out[24]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_25(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][25][0],w[0][25][1],w[0][25][2],w[0][25][3],w[0][25][4],w[0][25][5],w[0][25][6],w[0][25][7],w[0][25][8],w[0][25][9],w[0][25][10],w[0][25][11],w[0][25][12],w[0][25][13],w[0][25][14],w[0][25][15],w[0][25][16],w[0][25][17],w[0][25][18],w[0][25][19],w[0][25][20],w[0][25][21],w[0][25][22],w[0][25][23],w[0][25][24],w[0][25][25],w[0][25][26],w[0][25][27],w[0][25][28],w[0][25][29],w[0][25][30],w[0][25][31],b[0][25],out[25]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_26(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][26][0],w[0][26][1],w[0][26][2],w[0][26][3],w[0][26][4],w[0][26][5],w[0][26][6],w[0][26][7],w[0][26][8],w[0][26][9],w[0][26][10],w[0][26][11],w[0][26][12],w[0][26][13],w[0][26][14],w[0][26][15],w[0][26][16],w[0][26][17],w[0][26][18],w[0][26][19],w[0][26][20],w[0][26][21],w[0][26][22],w[0][26][23],w[0][26][24],w[0][26][25],w[0][26][26],w[0][26][27],w[0][26][28],w[0][26][29],w[0][26][30],w[0][26][31],b[0][26],out[26]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_27(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][27][0],w[0][27][1],w[0][27][2],w[0][27][3],w[0][27][4],w[0][27][5],w[0][27][6],w[0][27][7],w[0][27][8],w[0][27][9],w[0][27][10],w[0][27][11],w[0][27][12],w[0][27][13],w[0][27][14],w[0][27][15],w[0][27][16],w[0][27][17],w[0][27][18],w[0][27][19],w[0][27][20],w[0][27][21],w[0][27][22],w[0][27][23],w[0][27][24],w[0][27][25],w[0][27][26],w[0][27][27],w[0][27][28],w[0][27][29],w[0][27][30],w[0][27][31],b[0][27],out[27]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_28(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][28][0],w[0][28][1],w[0][28][2],w[0][28][3],w[0][28][4],w[0][28][5],w[0][28][6],w[0][28][7],w[0][28][8],w[0][28][9],w[0][28][10],w[0][28][11],w[0][28][12],w[0][28][13],w[0][28][14],w[0][28][15],w[0][28][16],w[0][28][17],w[0][28][18],w[0][28][19],w[0][28][20],w[0][28][21],w[0][28][22],w[0][28][23],w[0][28][24],w[0][28][25],w[0][28][26],w[0][28][27],w[0][28][28],w[0][28][29],w[0][28][30],w[0][28][31],b[0][28],out[28]);
neuron32 #(.sizein(sizein),.sizew(sizew),.sizeout(sizeout)) n0_29(relu,in[0],in[1],in[2],in[3],in[4],in[5],in[6],in[7],in[8],in[9],in[10],in[11],in[12],in[13],in[14],in[15],in[16],in[17],in[18],in[19],in[20],in[21],in[22],in[23],in[24],in[25],in[26],in[27],in[28],in[29],in[30],in[31],w[0][29][0],w[0][29][1],w[0][29][2],w[0][29][3],w[0][29][4],w[0][29][5],w[0][29][6],w[0][29][7],w[0][29][8],w[0][29][9],w[0][29][10],w[0][29][11],w[0][29][12],w[0][29][13],w[0][29][14],w[0][29][15],w[0][29][16],w[0][29][17],w[0][29][18],w[0][29][19],w[0][29][20],w[0][29][21],w[0][29][22],w[0][29][23],w[0][29][24],w[0][29][25],w[0][29][26],w[0][29][27],w[0][29][28],w[0][29][29],w[0][29][30],w[0][29][31],b[0][29],out[29]);

parameter IDLE=0;
parameter LOADIN=1;
parameter LOADIN0=2;
parameter LOADIN1=3;
parameter LOADW=4;
parameter LOADW0=5;
parameter LOADW1=6;
parameter LOADB=7;
parameter LOADB0=8;
parameter LOADB1=9;
parameter INIT=10;
parameter WAIT0=11;
parameter TRANS=12;
parameter WAIT1=13;
parameter RESULT=14;
parameter FINISH=15;

reg[7:0] state,prev_state;
reg[7:0] cin,cl,cn,cw;

reg[7:0] i;
reg[7:0] delay;

reg[sizeout-1:0] max;
reg[7:0] count,maxc;

assign debug=state;
assign debug1=w[0][2][3]|(b[0][5]<<8)|(w[1][4][5]<<16)|(b[1][6]<<24);

always@(posedge clk)begin
	if(rst)begin
		state<=IDLE;
	end
	else begin
		case(state)
		IDLE:begin
			if(start)begin
				cin<=0;
				cl<=0;
				cn<=0;
				cw<=0;
				relu<=1;
				finished<=0;
				state<=LOADIN;
			end
			else begin
				state<=IDLE;
			end
		end
		LOADIN:begin
			if(cin<32)begin
				rmode<=0;
				rs<=1;
				rin<=cin;
				state<=LOADIN0;
			end
			else begin
				cl<=1;
				cn<=0;
				cw<=0;
				rmode<=1;
				state<=LOADW;
			end
		end
		LOADIN0:begin
			rs<=0;
			state<=LOADIN1;
		end
		LOADIN1:begin
			if(rf)begin
				in[cin]<=ram_in;
				cin<=cin+1;
				state<=LOADIN;
			end
			else begin
				state<=LOADIN1;
			end
		end
		LOADW:begin
			if(cl==2)begin
				if(cn==10)begin
					cl<=2;
					cn<=0;
					cw<=0;
					rmode<=1;
					state<=LOADB;
				end
				else begin
					if(cw==32)begin
						cn<=cn+1;
						cw<=0;
						state<=LOADW;
					end
					else if(cw>=30)begin
						w[0][cn][cw]<=0;
						cw<=cw+1;
						state<=LOADW;
					end
					else begin
						rmode<=1;
						rs<=1;
						rlayer<=cl;
						rn<=cn;
						rin<=cw+1;
						cw<=cw+1;
						state<=LOADW0;
					end
				end
			end
			else if(cl==1)begin
				if(cn==30)begin
					//cl<=cl+1;
					cl<=1;
					cn<=0;
					cw<=0;
					rmode<=1;
					state<=LOADB;
				end
				else begin
					if(cw==32)begin
						cn<=cn+1;
						cw<=0;
						state<=LOADW;
					end
					else begin
						rmode<=1;
						rs<=1;
						rlayer<=cl;
						rn<=cn;
						rin<=cw+1;
						cw<=cw+1;
						state<=LOADW0;
					end
				end
			end
			else begin
				cl<=cl+1;
				state<=LOADW;
			end
		end
		LOADW0:begin
			rs<=0;
			state<=LOADW1;
		end
		LOADW1:begin
			if(rf)begin
				w[0][cn][cw-1]<=ram_w;
				state<=LOADW;
			end
			else begin
				state<=LOADW1;
			end
		end
		LOADB:begin
			if(cl==2)begin
				if(cn==10)begin
					cn<=0;
					cw<=0;
					delay<=10;
					state<=WAIT1;
				end
				else begin
					rmode<=1;
					rs<=1;
					rlayer<=cl;
					rn<=cn;
					rin<=0;
					cn<=cn+1;
					state<=LOADB0;
				end
			end
			else if(cl==1)begin
				if(cn==30)begin
					//cl<=cl+1;
					cn<=0;
					cw<=0;
					delay<=10;
					state<=WAIT0;
				end
				else begin
					rmode<=1;
					rs<=1;
					rlayer<=cl;
					rn<=cn;
					rin<=0;
					cn<=cn+1;
					state<=LOADB0;
				end
			end
			else begin
				cl<=cl+1;
				state<=LOADB;
			end
		end
		LOADB0:begin
			rs<=0;
			state<=LOADB1;
		end
		LOADB1:begin
			if(rf)begin
				b[0][cn-1]<=ram_w;
				state<=LOADB;
			end
			else begin
				state<=LOADB1;
			end
		end
		WAIT0:begin
			if(delay>0)begin
				delay<=delay-1;
			end
			else begin
				max<=0;
				count<=0;
				maxc<=0;
				cn<=0;
				state<=TRANS;
			end
		end
		TRANS:begin
			if(cn<30)begin
				outtemp[cn]<=out[cn];
				cn<=cn+1;
				state<=TRANS;
			end
			else if(cn<62)begin
				if(cn<60)begin
					in[cn-30]<=outtemp[cn-30];
				end
				else begin
					in[cn-30]<=0;
				end
				cn<=cn+1;
				state<=TRANS;
			end
			else begin
				cl<=2;
				rmode<=1;
				cn<=0;
				cw<=0;
				relu<=0;
				state<=LOADW;
			end
		end
		WAIT1:begin
			if(delay>0)begin
				delay<=delay-1;
			end
			else begin
				max<=0;
				count<=0;
				maxc<=0;
				state<=RESULT;
			end
		end
		RESULT:begin
			if(count<10)begin
				if(out[count][sizeout-1]==0)begin
					if(out[count][sizeout-2:0]>max)begin
						maxc<=count;
						max<=out[count][sizeout-2:0];
					end
				end
				count<=count+1;
				state<=RESULT;
			end
			else begin
				result<=maxc;
				state<=FINISH;
			end
		end
		FINISH:begin
			finished<=1;
			state<=IDLE;
		end
		endcase
	end
end

endmodule
